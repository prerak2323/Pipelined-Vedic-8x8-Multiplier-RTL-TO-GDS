module vedic8x8 (clk,
    ground,
    overflow,
    a,
    b,
    prod);
 input clk;
 input ground;
 output overflow;
 input [7:0] a;
 input [7:0] b;
 output [15:0] prod;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire c1;
 wire c1_s1;
 wire c1_s2;
 wire c2;
 wire c2_s2;
 wire ov1;
 wire ov2;
 wire ov3;
 wire ov4;
 wire \M0/c1 ;
 wire \M0/c2 ;
 wire \M0/cnet ;
 wire \M0/M0/a0b1 ;
 wire \M0/M0/a1b0 ;
 wire \M0/M0/a1b1 ;
 wire \M0/M0/carry ;
 wire \M0/M1/a0b1 ;
 wire \M0/M1/a1b0 ;
 wire \M0/M1/a1b1 ;
 wire \M0/M1/carry ;
 wire \M0/M2/a0b1 ;
 wire \M0/M2/a1b0 ;
 wire \M0/M2/a1b1 ;
 wire \M0/M2/carry ;
 wire \M0/M3/a0b1 ;
 wire \M0/M3/a1b0 ;
 wire \M0/M3/a1b1 ;
 wire \M0/M3/carry ;
 wire \M0/stage1/_00_ ;
 wire \M0/stage1/_01_ ;
 wire \M0/stage1/_02_ ;
 wire \M0/stage1/_03_ ;
 wire \M0/stage1/FA1_0/ha1_carry ;
 wire \M0/stage1/FA1_0/ha1_sum ;
 wire \M0/stage1/FA1_0/ha2_carry ;
 wire \M0/stage1/gen_csa[1].FA0/ha1_carry ;
 wire \M0/stage1/gen_csa[1].FA0/ha1_sum ;
 wire \M0/stage1/gen_csa[1].FA0/ha2_carry ;
 wire \M0/stage1/gen_csa[1].FA1/ha1_carry ;
 wire \M0/stage1/gen_csa[1].FA1/ha1_sum ;
 wire \M0/stage1/gen_csa[1].FA1/ha2_carry ;
 wire \M0/stage1/gen_csa[2].FA0/ha1_carry ;
 wire \M0/stage1/gen_csa[2].FA0/ha1_sum ;
 wire \M0/stage1/gen_csa[2].FA0/ha2_carry ;
 wire \M0/stage1/gen_csa[2].FA1/ha1_carry ;
 wire \M0/stage1/gen_csa[2].FA1/ha1_sum ;
 wire \M0/stage1/gen_csa[2].FA1/ha2_carry ;
 wire \M0/stage1/gen_csa[3].FA0/ha1_carry ;
 wire \M0/stage1/gen_csa[3].FA0/ha1_sum ;
 wire \M0/stage1/gen_csa[3].FA0/ha2_carry ;
 wire \M0/stage1/gen_csa[3].FA1/ha1_carry ;
 wire \M0/stage1/gen_csa[3].FA1/ha1_sum ;
 wire \M0/stage1/gen_csa[3].FA1/ha2_carry ;
 wire \M0/stage2/_00_ ;
 wire \M0/stage2/_01_ ;
 wire \M0/stage2/_02_ ;
 wire \M0/stage2/_03_ ;
 wire \M0/stage2/FA1_0/ha1_carry ;
 wire \M0/stage2/FA1_0/ha1_sum ;
 wire \M0/stage2/FA1_0/ha2_carry ;
 wire \M0/stage2/gen_csa[1].FA0/ha1_carry ;
 wire \M0/stage2/gen_csa[1].FA0/ha1_sum ;
 wire \M0/stage2/gen_csa[1].FA0/ha2_carry ;
 wire \M0/stage2/gen_csa[1].FA1/ha1_carry ;
 wire \M0/stage2/gen_csa[1].FA1/ha1_sum ;
 wire \M0/stage2/gen_csa[1].FA1/ha2_carry ;
 wire \M0/stage2/gen_csa[2].FA0/ha1_carry ;
 wire \M0/stage2/gen_csa[2].FA0/ha1_sum ;
 wire \M0/stage2/gen_csa[2].FA0/ha2_carry ;
 wire \M0/stage2/gen_csa[2].FA1/ha1_carry ;
 wire \M0/stage2/gen_csa[2].FA1/ha1_sum ;
 wire \M0/stage2/gen_csa[2].FA1/ha2_carry ;
 wire \M0/stage2/gen_csa[3].FA0/ha1_carry ;
 wire \M0/stage2/gen_csa[3].FA0/ha1_sum ;
 wire \M0/stage2/gen_csa[3].FA0/ha2_carry ;
 wire \M0/stage2/gen_csa[3].FA1/ha1_carry ;
 wire \M0/stage2/gen_csa[3].FA1/ha1_sum ;
 wire \M0/stage2/gen_csa[3].FA1/ha2_carry ;
 wire \M0/stage3/_00_ ;
 wire \M0/stage3/_01_ ;
 wire \M0/stage3/_02_ ;
 wire \M0/stage3/_03_ ;
 wire \M0/stage3/FA1_0/ha1_carry ;
 wire \M0/stage3/FA1_0/ha1_sum ;
 wire \M0/stage3/FA1_0/ha2_carry ;
 wire \M0/stage3/gen_csa[1].FA0/ha1_carry ;
 wire \M0/stage3/gen_csa[1].FA0/ha1_sum ;
 wire \M0/stage3/gen_csa[1].FA0/ha2_carry ;
 wire \M0/stage3/gen_csa[1].FA1/ha1_carry ;
 wire \M0/stage3/gen_csa[1].FA1/ha1_sum ;
 wire \M0/stage3/gen_csa[1].FA1/ha2_carry ;
 wire \M0/stage3/gen_csa[2].FA0/ha1_carry ;
 wire \M0/stage3/gen_csa[2].FA0/ha1_sum ;
 wire \M0/stage3/gen_csa[2].FA0/ha2_carry ;
 wire \M0/stage3/gen_csa[2].FA1/ha1_carry ;
 wire \M0/stage3/gen_csa[2].FA1/ha1_sum ;
 wire \M0/stage3/gen_csa[2].FA1/ha2_carry ;
 wire \M0/stage3/gen_csa[3].FA0/ha1_carry ;
 wire \M0/stage3/gen_csa[3].FA0/ha1_sum ;
 wire \M0/stage3/gen_csa[3].FA0/ha2_carry ;
 wire \M0/stage3/gen_csa[3].FA1/ha1_carry ;
 wire \M0/stage3/gen_csa[3].FA1/ha1_sum ;
 wire \M0/stage3/gen_csa[3].FA1/ha2_carry ;
 wire \M1/c1 ;
 wire \M1/c2 ;
 wire \M1/cnet ;
 wire \M1/M0/a0b1 ;
 wire \M1/M0/a1b0 ;
 wire \M1/M0/a1b1 ;
 wire \M1/M0/carry ;
 wire \M1/M1/a0b1 ;
 wire \M1/M1/a1b0 ;
 wire \M1/M1/a1b1 ;
 wire \M1/M1/carry ;
 wire \M1/M2/a0b1 ;
 wire \M1/M2/a1b0 ;
 wire \M1/M2/a1b1 ;
 wire \M1/M2/carry ;
 wire \M1/M3/a0b1 ;
 wire \M1/M3/a1b0 ;
 wire \M1/M3/a1b1 ;
 wire \M1/M3/carry ;
 wire \M1/stage1/_00_ ;
 wire \M1/stage1/_01_ ;
 wire \M1/stage1/_02_ ;
 wire \M1/stage1/_03_ ;
 wire \M1/stage1/FA1_0/ha1_carry ;
 wire \M1/stage1/FA1_0/ha1_sum ;
 wire \M1/stage1/FA1_0/ha2_carry ;
 wire \M1/stage1/gen_csa[1].FA0/ha1_carry ;
 wire \M1/stage1/gen_csa[1].FA0/ha1_sum ;
 wire \M1/stage1/gen_csa[1].FA0/ha2_carry ;
 wire \M1/stage1/gen_csa[1].FA1/ha1_carry ;
 wire \M1/stage1/gen_csa[1].FA1/ha1_sum ;
 wire \M1/stage1/gen_csa[1].FA1/ha2_carry ;
 wire \M1/stage1/gen_csa[2].FA0/ha1_carry ;
 wire \M1/stage1/gen_csa[2].FA0/ha1_sum ;
 wire \M1/stage1/gen_csa[2].FA0/ha2_carry ;
 wire \M1/stage1/gen_csa[2].FA1/ha1_carry ;
 wire \M1/stage1/gen_csa[2].FA1/ha1_sum ;
 wire \M1/stage1/gen_csa[2].FA1/ha2_carry ;
 wire \M1/stage1/gen_csa[3].FA0/ha1_carry ;
 wire \M1/stage1/gen_csa[3].FA0/ha1_sum ;
 wire \M1/stage1/gen_csa[3].FA0/ha2_carry ;
 wire \M1/stage1/gen_csa[3].FA1/ha1_carry ;
 wire \M1/stage1/gen_csa[3].FA1/ha1_sum ;
 wire \M1/stage1/gen_csa[3].FA1/ha2_carry ;
 wire \M1/stage2/_00_ ;
 wire \M1/stage2/_01_ ;
 wire \M1/stage2/_02_ ;
 wire \M1/stage2/_03_ ;
 wire \M1/stage2/FA1_0/ha1_carry ;
 wire \M1/stage2/FA1_0/ha1_sum ;
 wire \M1/stage2/FA1_0/ha2_carry ;
 wire \M1/stage2/gen_csa[1].FA0/ha1_carry ;
 wire \M1/stage2/gen_csa[1].FA0/ha1_sum ;
 wire \M1/stage2/gen_csa[1].FA0/ha2_carry ;
 wire \M1/stage2/gen_csa[1].FA1/ha1_carry ;
 wire \M1/stage2/gen_csa[1].FA1/ha1_sum ;
 wire \M1/stage2/gen_csa[1].FA1/ha2_carry ;
 wire \M1/stage2/gen_csa[2].FA0/ha1_carry ;
 wire \M1/stage2/gen_csa[2].FA0/ha1_sum ;
 wire \M1/stage2/gen_csa[2].FA0/ha2_carry ;
 wire \M1/stage2/gen_csa[2].FA1/ha1_carry ;
 wire \M1/stage2/gen_csa[2].FA1/ha1_sum ;
 wire \M1/stage2/gen_csa[2].FA1/ha2_carry ;
 wire \M1/stage2/gen_csa[3].FA0/ha1_carry ;
 wire \M1/stage2/gen_csa[3].FA0/ha1_sum ;
 wire \M1/stage2/gen_csa[3].FA0/ha2_carry ;
 wire \M1/stage2/gen_csa[3].FA1/ha1_carry ;
 wire \M1/stage2/gen_csa[3].FA1/ha1_sum ;
 wire \M1/stage2/gen_csa[3].FA1/ha2_carry ;
 wire \M1/stage3/_00_ ;
 wire \M1/stage3/_01_ ;
 wire \M1/stage3/_02_ ;
 wire \M1/stage3/_03_ ;
 wire \M1/stage3/FA1_0/ha1_carry ;
 wire \M1/stage3/FA1_0/ha1_sum ;
 wire \M1/stage3/FA1_0/ha2_carry ;
 wire \M1/stage3/gen_csa[1].FA0/ha1_carry ;
 wire \M1/stage3/gen_csa[1].FA0/ha1_sum ;
 wire \M1/stage3/gen_csa[1].FA0/ha2_carry ;
 wire \M1/stage3/gen_csa[1].FA1/ha1_carry ;
 wire \M1/stage3/gen_csa[1].FA1/ha1_sum ;
 wire \M1/stage3/gen_csa[1].FA1/ha2_carry ;
 wire \M1/stage3/gen_csa[2].FA0/ha1_carry ;
 wire \M1/stage3/gen_csa[2].FA0/ha1_sum ;
 wire \M1/stage3/gen_csa[2].FA0/ha2_carry ;
 wire \M1/stage3/gen_csa[2].FA1/ha1_carry ;
 wire \M1/stage3/gen_csa[2].FA1/ha1_sum ;
 wire \M1/stage3/gen_csa[2].FA1/ha2_carry ;
 wire \M1/stage3/gen_csa[3].FA0/ha1_carry ;
 wire \M1/stage3/gen_csa[3].FA0/ha1_sum ;
 wire \M1/stage3/gen_csa[3].FA0/ha2_carry ;
 wire \M1/stage3/gen_csa[3].FA1/ha1_carry ;
 wire \M1/stage3/gen_csa[3].FA1/ha1_sum ;
 wire \M1/stage3/gen_csa[3].FA1/ha2_carry ;
 wire \M2/c1 ;
 wire \M2/c2 ;
 wire \M2/cnet ;
 wire \M2/M0/a0b1 ;
 wire \M2/M0/a1b0 ;
 wire \M2/M0/a1b1 ;
 wire \M2/M0/carry ;
 wire \M2/M1/a0b1 ;
 wire \M2/M1/a1b0 ;
 wire \M2/M1/a1b1 ;
 wire \M2/M1/carry ;
 wire \M2/M2/a0b1 ;
 wire \M2/M2/a1b0 ;
 wire \M2/M2/a1b1 ;
 wire \M2/M2/carry ;
 wire \M2/M3/a0b1 ;
 wire \M2/M3/a1b0 ;
 wire \M2/M3/a1b1 ;
 wire \M2/M3/carry ;
 wire \M2/stage1/_00_ ;
 wire \M2/stage1/_01_ ;
 wire \M2/stage1/_02_ ;
 wire \M2/stage1/_03_ ;
 wire \M2/stage1/FA1_0/ha1_carry ;
 wire \M2/stage1/FA1_0/ha1_sum ;
 wire \M2/stage1/FA1_0/ha2_carry ;
 wire \M2/stage1/gen_csa[1].FA0/ha1_carry ;
 wire \M2/stage1/gen_csa[1].FA0/ha1_sum ;
 wire \M2/stage1/gen_csa[1].FA0/ha2_carry ;
 wire \M2/stage1/gen_csa[1].FA1/ha1_carry ;
 wire \M2/stage1/gen_csa[1].FA1/ha1_sum ;
 wire \M2/stage1/gen_csa[1].FA1/ha2_carry ;
 wire \M2/stage1/gen_csa[2].FA0/ha1_carry ;
 wire \M2/stage1/gen_csa[2].FA0/ha1_sum ;
 wire \M2/stage1/gen_csa[2].FA0/ha2_carry ;
 wire \M2/stage1/gen_csa[2].FA1/ha1_carry ;
 wire \M2/stage1/gen_csa[2].FA1/ha1_sum ;
 wire \M2/stage1/gen_csa[2].FA1/ha2_carry ;
 wire \M2/stage1/gen_csa[3].FA0/ha1_carry ;
 wire \M2/stage1/gen_csa[3].FA0/ha1_sum ;
 wire \M2/stage1/gen_csa[3].FA0/ha2_carry ;
 wire \M2/stage1/gen_csa[3].FA1/ha1_carry ;
 wire \M2/stage1/gen_csa[3].FA1/ha1_sum ;
 wire \M2/stage1/gen_csa[3].FA1/ha2_carry ;
 wire \M2/stage2/_00_ ;
 wire \M2/stage2/_01_ ;
 wire \M2/stage2/_02_ ;
 wire \M2/stage2/_03_ ;
 wire \M2/stage2/FA1_0/ha1_carry ;
 wire \M2/stage2/FA1_0/ha1_sum ;
 wire \M2/stage2/FA1_0/ha2_carry ;
 wire \M2/stage2/gen_csa[1].FA0/ha1_carry ;
 wire \M2/stage2/gen_csa[1].FA0/ha1_sum ;
 wire \M2/stage2/gen_csa[1].FA0/ha2_carry ;
 wire \M2/stage2/gen_csa[1].FA1/ha1_carry ;
 wire \M2/stage2/gen_csa[1].FA1/ha1_sum ;
 wire \M2/stage2/gen_csa[1].FA1/ha2_carry ;
 wire \M2/stage2/gen_csa[2].FA0/ha1_carry ;
 wire \M2/stage2/gen_csa[2].FA0/ha1_sum ;
 wire \M2/stage2/gen_csa[2].FA0/ha2_carry ;
 wire \M2/stage2/gen_csa[2].FA1/ha1_carry ;
 wire \M2/stage2/gen_csa[2].FA1/ha1_sum ;
 wire \M2/stage2/gen_csa[2].FA1/ha2_carry ;
 wire \M2/stage2/gen_csa[3].FA0/ha1_carry ;
 wire \M2/stage2/gen_csa[3].FA0/ha1_sum ;
 wire \M2/stage2/gen_csa[3].FA0/ha2_carry ;
 wire \M2/stage2/gen_csa[3].FA1/ha1_carry ;
 wire \M2/stage2/gen_csa[3].FA1/ha1_sum ;
 wire \M2/stage2/gen_csa[3].FA1/ha2_carry ;
 wire \M2/stage3/_00_ ;
 wire \M2/stage3/_01_ ;
 wire \M2/stage3/_02_ ;
 wire \M2/stage3/_03_ ;
 wire \M2/stage3/FA1_0/ha1_carry ;
 wire \M2/stage3/FA1_0/ha1_sum ;
 wire \M2/stage3/FA1_0/ha2_carry ;
 wire \M2/stage3/gen_csa[1].FA0/ha1_carry ;
 wire \M2/stage3/gen_csa[1].FA0/ha1_sum ;
 wire \M2/stage3/gen_csa[1].FA0/ha2_carry ;
 wire \M2/stage3/gen_csa[1].FA1/ha1_carry ;
 wire \M2/stage3/gen_csa[1].FA1/ha1_sum ;
 wire \M2/stage3/gen_csa[1].FA1/ha2_carry ;
 wire \M2/stage3/gen_csa[2].FA0/ha1_carry ;
 wire \M2/stage3/gen_csa[2].FA0/ha1_sum ;
 wire \M2/stage3/gen_csa[2].FA0/ha2_carry ;
 wire \M2/stage3/gen_csa[2].FA1/ha1_carry ;
 wire \M2/stage3/gen_csa[2].FA1/ha1_sum ;
 wire \M2/stage3/gen_csa[2].FA1/ha2_carry ;
 wire \M2/stage3/gen_csa[3].FA0/ha1_carry ;
 wire \M2/stage3/gen_csa[3].FA0/ha1_sum ;
 wire \M2/stage3/gen_csa[3].FA0/ha2_carry ;
 wire \M2/stage3/gen_csa[3].FA1/ha1_carry ;
 wire \M2/stage3/gen_csa[3].FA1/ha1_sum ;
 wire \M2/stage3/gen_csa[3].FA1/ha2_carry ;
 wire \M3/c1 ;
 wire \M3/c2 ;
 wire \M3/cnet ;
 wire \M3/M0/a0b1 ;
 wire \M3/M0/a1b0 ;
 wire \M3/M0/a1b1 ;
 wire \M3/M0/carry ;
 wire \M3/M1/a0b1 ;
 wire \M3/M1/a1b0 ;
 wire \M3/M1/a1b1 ;
 wire \M3/M1/carry ;
 wire \M3/M2/a0b1 ;
 wire \M3/M2/a1b0 ;
 wire \M3/M2/a1b1 ;
 wire \M3/M2/carry ;
 wire \M3/M3/a0b1 ;
 wire \M3/M3/a1b0 ;
 wire \M3/M3/a1b1 ;
 wire \M3/M3/carry ;
 wire \M3/stage1/_00_ ;
 wire \M3/stage1/_01_ ;
 wire \M3/stage1/_02_ ;
 wire \M3/stage1/_03_ ;
 wire \M3/stage1/FA1_0/ha1_carry ;
 wire \M3/stage1/FA1_0/ha1_sum ;
 wire \M3/stage1/FA1_0/ha2_carry ;
 wire \M3/stage1/gen_csa[1].FA0/ha1_carry ;
 wire \M3/stage1/gen_csa[1].FA0/ha1_sum ;
 wire \M3/stage1/gen_csa[1].FA0/ha2_carry ;
 wire \M3/stage1/gen_csa[1].FA1/ha1_carry ;
 wire \M3/stage1/gen_csa[1].FA1/ha1_sum ;
 wire \M3/stage1/gen_csa[1].FA1/ha2_carry ;
 wire \M3/stage1/gen_csa[2].FA0/ha1_carry ;
 wire \M3/stage1/gen_csa[2].FA0/ha1_sum ;
 wire \M3/stage1/gen_csa[2].FA0/ha2_carry ;
 wire \M3/stage1/gen_csa[2].FA1/ha1_carry ;
 wire \M3/stage1/gen_csa[2].FA1/ha1_sum ;
 wire \M3/stage1/gen_csa[2].FA1/ha2_carry ;
 wire \M3/stage1/gen_csa[3].FA0/ha1_carry ;
 wire \M3/stage1/gen_csa[3].FA0/ha1_sum ;
 wire \M3/stage1/gen_csa[3].FA0/ha2_carry ;
 wire \M3/stage1/gen_csa[3].FA1/ha1_carry ;
 wire \M3/stage1/gen_csa[3].FA1/ha1_sum ;
 wire \M3/stage1/gen_csa[3].FA1/ha2_carry ;
 wire \M3/stage2/_00_ ;
 wire \M3/stage2/_01_ ;
 wire \M3/stage2/_02_ ;
 wire \M3/stage2/_03_ ;
 wire \M3/stage2/FA1_0/ha1_carry ;
 wire \M3/stage2/FA1_0/ha1_sum ;
 wire \M3/stage2/FA1_0/ha2_carry ;
 wire \M3/stage2/gen_csa[1].FA0/ha1_carry ;
 wire \M3/stage2/gen_csa[1].FA0/ha1_sum ;
 wire \M3/stage2/gen_csa[1].FA0/ha2_carry ;
 wire \M3/stage2/gen_csa[1].FA1/ha1_carry ;
 wire \M3/stage2/gen_csa[1].FA1/ha1_sum ;
 wire \M3/stage2/gen_csa[1].FA1/ha2_carry ;
 wire \M3/stage2/gen_csa[2].FA0/ha1_carry ;
 wire \M3/stage2/gen_csa[2].FA0/ha1_sum ;
 wire \M3/stage2/gen_csa[2].FA0/ha2_carry ;
 wire \M3/stage2/gen_csa[2].FA1/ha1_carry ;
 wire \M3/stage2/gen_csa[2].FA1/ha1_sum ;
 wire \M3/stage2/gen_csa[2].FA1/ha2_carry ;
 wire \M3/stage2/gen_csa[3].FA0/ha1_carry ;
 wire \M3/stage2/gen_csa[3].FA0/ha1_sum ;
 wire \M3/stage2/gen_csa[3].FA0/ha2_carry ;
 wire \M3/stage2/gen_csa[3].FA1/ha1_carry ;
 wire \M3/stage2/gen_csa[3].FA1/ha1_sum ;
 wire \M3/stage2/gen_csa[3].FA1/ha2_carry ;
 wire \M3/stage3/_00_ ;
 wire \M3/stage3/_01_ ;
 wire \M3/stage3/_02_ ;
 wire \M3/stage3/_03_ ;
 wire \M3/stage3/FA1_0/ha1_carry ;
 wire \M3/stage3/FA1_0/ha1_sum ;
 wire \M3/stage3/FA1_0/ha2_carry ;
 wire \M3/stage3/gen_csa[1].FA0/ha1_carry ;
 wire \M3/stage3/gen_csa[1].FA0/ha1_sum ;
 wire \M3/stage3/gen_csa[1].FA0/ha2_carry ;
 wire \M3/stage3/gen_csa[1].FA1/ha1_carry ;
 wire \M3/stage3/gen_csa[1].FA1/ha1_sum ;
 wire \M3/stage3/gen_csa[1].FA1/ha2_carry ;
 wire \M3/stage3/gen_csa[2].FA0/ha1_carry ;
 wire \M3/stage3/gen_csa[2].FA0/ha1_sum ;
 wire \M3/stage3/gen_csa[2].FA0/ha2_carry ;
 wire \M3/stage3/gen_csa[2].FA1/ha1_carry ;
 wire \M3/stage3/gen_csa[2].FA1/ha1_sum ;
 wire \M3/stage3/gen_csa[2].FA1/ha2_carry ;
 wire \M3/stage3/gen_csa[3].FA0/ha1_carry ;
 wire \M3/stage3/gen_csa[3].FA0/ha1_sum ;
 wire \M3/stage3/gen_csa[3].FA0/ha2_carry ;
 wire \M3/stage3/gen_csa[3].FA1/ha1_carry ;
 wire \M3/stage3/gen_csa[3].FA1/ha1_sum ;
 wire \M3/stage3/gen_csa[3].FA1/ha2_carry ;
 wire \stage1/_00_ ;
 wire \stage1/_01_ ;
 wire \stage1/_02_ ;
 wire \stage1/_03_ ;
 wire \stage1/_04_ ;
 wire \stage1/_05_ ;
 wire \stage1/_06_ ;
 wire \stage1/_07_ ;
 wire \stage1/FA1_0/ha1_carry ;
 wire \stage1/FA1_0/ha1_sum ;
 wire \stage1/FA1_0/ha2_carry ;
 wire \stage1/gen_csa[1].FA0/ha1_carry ;
 wire \stage1/gen_csa[1].FA0/ha1_sum ;
 wire \stage1/gen_csa[1].FA0/ha2_carry ;
 wire \stage1/gen_csa[1].FA1/ha1_carry ;
 wire \stage1/gen_csa[1].FA1/ha1_sum ;
 wire \stage1/gen_csa[1].FA1/ha2_carry ;
 wire \stage1/gen_csa[2].FA0/ha1_carry ;
 wire \stage1/gen_csa[2].FA0/ha1_sum ;
 wire \stage1/gen_csa[2].FA0/ha2_carry ;
 wire \stage1/gen_csa[2].FA1/ha1_carry ;
 wire \stage1/gen_csa[2].FA1/ha1_sum ;
 wire \stage1/gen_csa[2].FA1/ha2_carry ;
 wire \stage1/gen_csa[3].FA0/ha1_carry ;
 wire \stage1/gen_csa[3].FA0/ha1_sum ;
 wire \stage1/gen_csa[3].FA0/ha2_carry ;
 wire \stage1/gen_csa[3].FA1/ha1_carry ;
 wire \stage1/gen_csa[3].FA1/ha1_sum ;
 wire \stage1/gen_csa[3].FA1/ha2_carry ;
 wire \stage1/gen_csa[4].FA0/ha1_carry ;
 wire \stage1/gen_csa[4].FA0/ha1_sum ;
 wire \stage1/gen_csa[4].FA0/ha2_carry ;
 wire \stage1/gen_csa[4].FA1/ha1_carry ;
 wire \stage1/gen_csa[4].FA1/ha1_sum ;
 wire \stage1/gen_csa[4].FA1/ha2_carry ;
 wire \stage1/gen_csa[5].FA0/ha1_carry ;
 wire \stage1/gen_csa[5].FA0/ha1_sum ;
 wire \stage1/gen_csa[5].FA0/ha2_carry ;
 wire \stage1/gen_csa[5].FA1/ha1_carry ;
 wire \stage1/gen_csa[5].FA1/ha1_sum ;
 wire \stage1/gen_csa[5].FA1/ha2_carry ;
 wire \stage1/gen_csa[6].FA0/ha1_carry ;
 wire \stage1/gen_csa[6].FA0/ha1_sum ;
 wire \stage1/gen_csa[6].FA0/ha2_carry ;
 wire \stage1/gen_csa[6].FA1/ha1_carry ;
 wire \stage1/gen_csa[6].FA1/ha1_sum ;
 wire \stage1/gen_csa[6].FA1/ha2_carry ;
 wire \stage1/gen_csa[7].FA0/ha1_carry ;
 wire \stage1/gen_csa[7].FA0/ha1_sum ;
 wire \stage1/gen_csa[7].FA0/ha2_carry ;
 wire \stage1/gen_csa[7].FA1/ha1_carry ;
 wire \stage1/gen_csa[7].FA1/ha1_sum ;
 wire \stage1/gen_csa[7].FA1/ha2_carry ;
 wire \stage2/_00_ ;
 wire \stage2/_01_ ;
 wire \stage2/_02_ ;
 wire \stage2/_03_ ;
 wire \stage2/_04_ ;
 wire \stage2/_05_ ;
 wire \stage2/_06_ ;
 wire \stage2/_07_ ;
 wire \stage2/FA1_0/ha1_carry ;
 wire \stage2/FA1_0/ha1_sum ;
 wire \stage2/FA1_0/ha2_carry ;
 wire \stage2/gen_csa[1].FA0/ha1_carry ;
 wire \stage2/gen_csa[1].FA0/ha1_sum ;
 wire \stage2/gen_csa[1].FA0/ha2_carry ;
 wire \stage2/gen_csa[1].FA1/ha1_carry ;
 wire \stage2/gen_csa[1].FA1/ha1_sum ;
 wire \stage2/gen_csa[1].FA1/ha2_carry ;
 wire \stage2/gen_csa[2].FA0/ha1_carry ;
 wire \stage2/gen_csa[2].FA0/ha1_sum ;
 wire \stage2/gen_csa[2].FA0/ha2_carry ;
 wire \stage2/gen_csa[2].FA1/ha1_carry ;
 wire \stage2/gen_csa[2].FA1/ha1_sum ;
 wire \stage2/gen_csa[2].FA1/ha2_carry ;
 wire \stage2/gen_csa[3].FA0/ha1_carry ;
 wire \stage2/gen_csa[3].FA0/ha1_sum ;
 wire \stage2/gen_csa[3].FA0/ha2_carry ;
 wire \stage2/gen_csa[3].FA1/ha1_carry ;
 wire \stage2/gen_csa[3].FA1/ha1_sum ;
 wire \stage2/gen_csa[3].FA1/ha2_carry ;
 wire \stage2/gen_csa[4].FA0/ha1_carry ;
 wire \stage2/gen_csa[4].FA0/ha1_sum ;
 wire \stage2/gen_csa[4].FA0/ha2_carry ;
 wire \stage2/gen_csa[4].FA1/ha1_carry ;
 wire \stage2/gen_csa[4].FA1/ha1_sum ;
 wire \stage2/gen_csa[4].FA1/ha2_carry ;
 wire \stage2/gen_csa[5].FA0/ha1_carry ;
 wire \stage2/gen_csa[5].FA0/ha1_sum ;
 wire \stage2/gen_csa[5].FA0/ha2_carry ;
 wire \stage2/gen_csa[5].FA1/ha1_carry ;
 wire \stage2/gen_csa[5].FA1/ha1_sum ;
 wire \stage2/gen_csa[5].FA1/ha2_carry ;
 wire \stage2/gen_csa[6].FA0/ha1_carry ;
 wire \stage2/gen_csa[6].FA0/ha1_sum ;
 wire \stage2/gen_csa[6].FA0/ha2_carry ;
 wire \stage2/gen_csa[6].FA1/ha1_carry ;
 wire \stage2/gen_csa[6].FA1/ha1_sum ;
 wire \stage2/gen_csa[6].FA1/ha2_carry ;
 wire \stage2/gen_csa[7].FA0/ha1_carry ;
 wire \stage2/gen_csa[7].FA0/ha1_sum ;
 wire \stage2/gen_csa[7].FA0/ha2_carry ;
 wire \stage2/gen_csa[7].FA1/ha1_carry ;
 wire \stage2/gen_csa[7].FA1/ha1_sum ;
 wire \stage2/gen_csa[7].FA1/ha2_carry ;
 wire \stage3/_00_ ;
 wire \stage3/_01_ ;
 wire \stage3/_02_ ;
 wire \stage3/_03_ ;
 wire \stage3/_04_ ;
 wire \stage3/_05_ ;
 wire \stage3/_06_ ;
 wire \stage3/_07_ ;
 wire \stage3/FA1_0/ha1_carry ;
 wire \stage3/FA1_0/ha1_sum ;
 wire \stage3/FA1_0/ha2_carry ;
 wire \stage3/gen_csa[1].FA0/ha1_carry ;
 wire \stage3/gen_csa[1].FA0/ha1_sum ;
 wire \stage3/gen_csa[1].FA0/ha2_carry ;
 wire \stage3/gen_csa[1].FA1/ha1_carry ;
 wire \stage3/gen_csa[1].FA1/ha1_sum ;
 wire \stage3/gen_csa[1].FA1/ha2_carry ;
 wire \stage3/gen_csa[2].FA0/ha1_carry ;
 wire \stage3/gen_csa[2].FA0/ha1_sum ;
 wire \stage3/gen_csa[2].FA0/ha2_carry ;
 wire \stage3/gen_csa[2].FA1/ha1_carry ;
 wire \stage3/gen_csa[2].FA1/ha1_sum ;
 wire \stage3/gen_csa[2].FA1/ha2_carry ;
 wire \stage3/gen_csa[3].FA0/ha1_carry ;
 wire \stage3/gen_csa[3].FA0/ha1_sum ;
 wire \stage3/gen_csa[3].FA0/ha2_carry ;
 wire \stage3/gen_csa[3].FA1/ha1_carry ;
 wire \stage3/gen_csa[3].FA1/ha1_sum ;
 wire \stage3/gen_csa[3].FA1/ha2_carry ;
 wire \stage3/gen_csa[4].FA0/ha1_carry ;
 wire \stage3/gen_csa[4].FA0/ha1_sum ;
 wire \stage3/gen_csa[4].FA0/ha2_carry ;
 wire \stage3/gen_csa[4].FA1/ha1_carry ;
 wire \stage3/gen_csa[4].FA1/ha1_sum ;
 wire \stage3/gen_csa[4].FA1/ha2_carry ;
 wire \stage3/gen_csa[5].FA0/ha1_carry ;
 wire \stage3/gen_csa[5].FA0/ha1_sum ;
 wire \stage3/gen_csa[5].FA0/ha2_carry ;
 wire \stage3/gen_csa[5].FA1/ha1_carry ;
 wire \stage3/gen_csa[5].FA1/ha1_sum ;
 wire \stage3/gen_csa[5].FA1/ha2_carry ;
 wire \stage3/gen_csa[6].FA0/ha1_carry ;
 wire \stage3/gen_csa[6].FA0/ha1_sum ;
 wire \stage3/gen_csa[6].FA0/ha2_carry ;
 wire \stage3/gen_csa[6].FA1/ha1_carry ;
 wire \stage3/gen_csa[6].FA1/ha1_sum ;
 wire \stage3/gen_csa[6].FA1/ha2_carry ;
 wire \stage3/gen_csa[7].FA0/ha1_carry ;
 wire \stage3/gen_csa[7].FA0/ha1_sum ;
 wire \stage3/gen_csa[7].FA0/ha2_carry ;
 wire \stage3/gen_csa[7].FA1/ha1_carry ;
 wire \stage3/gen_csa[7].FA1/ha1_sum ;
 wire \stage3/gen_csa[7].FA1/ha2_carry ;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire [3:0] \M0/prodm0 ;
 wire [3:0] \M0/prodm1 ;
 wire [3:0] \M0/prodm2 ;
 wire [3:0] \M0/prodm3 ;
 wire [3:0] \M0/stage1/carry0 ;
 wire [3:0] \M0/stage1/carry1 ;
 wire [3:0] \M0/stage1/sum0 ;
 wire [3:0] \M0/stage1/sum1 ;
 wire [3:0] \M0/stage2/carry0 ;
 wire [3:0] \M0/stage2/carry1 ;
 wire [3:0] \M0/stage2/sum0 ;
 wire [3:0] \M0/stage2/sum1 ;
 wire [3:0] \M0/stage3/carry0 ;
 wire [3:0] \M0/stage3/carry1 ;
 wire [3:0] \M0/stage3/sum0 ;
 wire [3:0] \M0/stage3/sum1 ;
 wire [3:0] \M0/sums1 ;
 wire [3:0] \M0/sums2 ;
 wire [3:0] \M1/prodm0 ;
 wire [3:0] \M1/prodm1 ;
 wire [3:0] \M1/prodm2 ;
 wire [3:0] \M1/prodm3 ;
 wire [3:0] \M1/stage1/carry0 ;
 wire [3:0] \M1/stage1/carry1 ;
 wire [3:0] \M1/stage1/sum0 ;
 wire [3:0] \M1/stage1/sum1 ;
 wire [3:0] \M1/stage2/carry0 ;
 wire [3:0] \M1/stage2/carry1 ;
 wire [3:0] \M1/stage2/sum0 ;
 wire [3:0] \M1/stage2/sum1 ;
 wire [3:0] \M1/stage3/carry0 ;
 wire [3:0] \M1/stage3/carry1 ;
 wire [3:0] \M1/stage3/sum0 ;
 wire [3:0] \M1/stage3/sum1 ;
 wire [3:0] \M1/sums1 ;
 wire [3:0] \M1/sums2 ;
 wire [3:0] \M2/prodm0 ;
 wire [3:0] \M2/prodm1 ;
 wire [3:0] \M2/prodm2 ;
 wire [3:0] \M2/prodm3 ;
 wire [3:0] \M2/stage1/carry0 ;
 wire [3:0] \M2/stage1/carry1 ;
 wire [3:0] \M2/stage1/sum0 ;
 wire [3:0] \M2/stage1/sum1 ;
 wire [3:0] \M2/stage2/carry0 ;
 wire [3:0] \M2/stage2/carry1 ;
 wire [3:0] \M2/stage2/sum0 ;
 wire [3:0] \M2/stage2/sum1 ;
 wire [3:0] \M2/stage3/carry0 ;
 wire [3:0] \M2/stage3/carry1 ;
 wire [3:0] \M2/stage3/sum0 ;
 wire [3:0] \M2/stage3/sum1 ;
 wire [3:0] \M2/sums1 ;
 wire [3:0] \M2/sums2 ;
 wire [3:0] \M3/prodm0 ;
 wire [3:0] \M3/prodm1 ;
 wire [3:0] \M3/prodm2 ;
 wire [3:0] \M3/prodm3 ;
 wire [3:0] \M3/stage1/carry0 ;
 wire [3:0] \M3/stage1/carry1 ;
 wire [3:0] \M3/stage1/sum0 ;
 wire [3:0] \M3/stage1/sum1 ;
 wire [3:0] \M3/stage2/carry0 ;
 wire [3:0] \M3/stage2/carry1 ;
 wire [3:0] \M3/stage2/sum0 ;
 wire [3:0] \M3/stage2/sum1 ;
 wire [3:0] \M3/stage3/carry0 ;
 wire [3:0] \M3/stage3/carry1 ;
 wire [3:0] \M3/stage3/sum0 ;
 wire [3:0] \M3/stage3/sum1 ;
 wire [3:0] \M3/sums1 ;
 wire [3:0] \M3/sums2 ;
 wire [7:0] prodm0;
 wire [7:0] prodm0_s0;
 wire [7:0] prodm0_s1;
 wire [7:0] prodm0_s2;
 wire [7:0] prodm1;
 wire [7:0] prodm1_s0;
 wire [7:0] prodm2;
 wire [7:0] prodm2_s0;
 wire [7:0] prodm3;
 wire [7:0] prodm3_s0;
 wire [7:0] prodm3_s1;
 wire [7:0] prodm3_s2;
 wire [7:0] \stage1/carry0 ;
 wire [7:0] \stage1/carry1 ;
 wire [7:0] \stage1/sum0 ;
 wire [7:0] \stage1/sum1 ;
 wire [7:0] \stage2/carry0 ;
 wire [7:0] \stage2/carry1 ;
 wire [7:0] \stage2/sum0 ;
 wire [7:0] \stage2/sum1 ;
 wire [7:0] \stage3/carry0 ;
 wire [7:0] \stage3/carry1 ;
 wire [7:0] \stage3/sum0 ;
 wire [7:0] \stage3/sum1 ;
 wire [7:0] sum_s1;
 wire [7:0] sum_s2;
 wire [7:0] sums1;
 wire [7:0] sums2;
 wire [7:0] sums3;

 AND2_X1 \M0/M0/HA0/_0_  (.A1(\M0/M0/a0b1 ),
    .A2(\M0/M0/a1b0 ),
    .ZN(\M0/M0/carry ));
 XOR2_X2 \M0/M0/HA0/_1_  (.A(\M0/M0/a0b1 ),
    .B(\M0/M0/a1b0 ),
    .Z(prodm0[1]));
 AND2_X1 \M0/M0/HA1/_0_  (.A1(\M0/M0/a1b1 ),
    .A2(\M0/M0/carry ),
    .ZN(\M0/prodm0 [3]));
 XOR2_X2 \M0/M0/HA1/_1_  (.A(\M0/M0/a1b1 ),
    .B(\M0/M0/carry ),
    .Z(\M0/prodm0 [2]));
 AND2_X1 \M0/M0/_0_  (.A1(a[1]),
    .A2(b[1]),
    .ZN(\M0/M0/a1b1 ));
 AND2_X1 \M0/M0/_1_  (.A1(b[1]),
    .A2(a[0]),
    .ZN(\M0/M0/a0b1 ));
 AND2_X1 \M0/M0/_2_  (.A1(a[1]),
    .A2(b[0]),
    .ZN(\M0/M0/a1b0 ));
 AND2_X1 \M0/M0/_3_  (.A1(a[0]),
    .A2(b[0]),
    .ZN(prodm0[0]));
 AND2_X1 \M0/M1/HA0/_0_  (.A1(\M0/M1/a0b1 ),
    .A2(\M0/M1/a1b0 ),
    .ZN(\M0/M1/carry ));
 XOR2_X2 \M0/M1/HA0/_1_  (.A(\M0/M1/a0b1 ),
    .B(\M0/M1/a1b0 ),
    .Z(\M0/prodm1 [1]));
 AND2_X1 \M0/M1/HA1/_0_  (.A1(\M0/M1/a1b1 ),
    .A2(\M0/M1/carry ),
    .ZN(\M0/prodm1 [3]));
 XOR2_X2 \M0/M1/HA1/_1_  (.A(\M0/M1/a1b1 ),
    .B(\M0/M1/carry ),
    .Z(\M0/prodm1 [2]));
 AND2_X1 \M0/M1/_0_  (.A1(a[1]),
    .A2(b[3]),
    .ZN(\M0/M1/a1b1 ));
 AND2_X1 \M0/M1/_1_  (.A1(b[3]),
    .A2(a[0]),
    .ZN(\M0/M1/a0b1 ));
 AND2_X1 \M0/M1/_2_  (.A1(a[1]),
    .A2(b[2]),
    .ZN(\M0/M1/a1b0 ));
 AND2_X1 \M0/M1/_3_  (.A1(a[0]),
    .A2(b[2]),
    .ZN(\M0/prodm1 [0]));
 AND2_X1 \M0/M2/HA0/_0_  (.A1(\M0/M2/a0b1 ),
    .A2(\M0/M2/a1b0 ),
    .ZN(\M0/M2/carry ));
 XOR2_X2 \M0/M2/HA0/_1_  (.A(\M0/M2/a0b1 ),
    .B(\M0/M2/a1b0 ),
    .Z(\M0/prodm2 [1]));
 AND2_X1 \M0/M2/HA1/_0_  (.A1(\M0/M2/a1b1 ),
    .A2(\M0/M2/carry ),
    .ZN(\M0/prodm2 [3]));
 XOR2_X2 \M0/M2/HA1/_1_  (.A(\M0/M2/a1b1 ),
    .B(\M0/M2/carry ),
    .Z(\M0/prodm2 [2]));
 AND2_X1 \M0/M2/_0_  (.A1(a[3]),
    .A2(b[1]),
    .ZN(\M0/M2/a1b1 ));
 AND2_X1 \M0/M2/_1_  (.A1(b[1]),
    .A2(a[2]),
    .ZN(\M0/M2/a0b1 ));
 AND2_X1 \M0/M2/_2_  (.A1(a[3]),
    .A2(b[0]),
    .ZN(\M0/M2/a1b0 ));
 AND2_X1 \M0/M2/_3_  (.A1(a[2]),
    .A2(b[0]),
    .ZN(\M0/prodm2 [0]));
 AND2_X1 \M0/M3/HA0/_0_  (.A1(\M0/M3/a0b1 ),
    .A2(\M0/M3/a1b0 ),
    .ZN(\M0/M3/carry ));
 XOR2_X2 \M0/M3/HA0/_1_  (.A(\M0/M3/a0b1 ),
    .B(\M0/M3/a1b0 ),
    .Z(\M0/prodm3 [1]));
 AND2_X1 \M0/M3/HA1/_0_  (.A1(\M0/M3/a1b1 ),
    .A2(\M0/M3/carry ),
    .ZN(\M0/prodm3 [3]));
 XOR2_X2 \M0/M3/HA1/_1_  (.A(\M0/M3/a1b1 ),
    .B(\M0/M3/carry ),
    .Z(\M0/prodm3 [2]));
 AND2_X1 \M0/M3/_0_  (.A1(a[3]),
    .A2(b[3]),
    .ZN(\M0/M3/a1b1 ));
 AND2_X1 \M0/M3/_1_  (.A1(b[3]),
    .A2(a[2]),
    .ZN(\M0/M3/a0b1 ));
 AND2_X1 \M0/M3/_2_  (.A1(a[3]),
    .A2(b[2]),
    .ZN(\M0/M3/a1b0 ));
 AND2_X1 \M0/M3/_3_  (.A1(a[2]),
    .A2(b[2]),
    .ZN(\M0/prodm3 [0]));
 OR2_X2 \M0/_0_  (.A1(\M0/c1 ),
    .A2(\M0/c2 ),
    .ZN(\M0/cnet ));
 AND2_X1 \M0/stage1/FA1_0/HA1/_0_  (.A1(\M0/prodm1 [0]),
    .A2(\M0/prodm2 [0]),
    .ZN(\M0/stage1/FA1_0/ha1_carry ));
 XOR2_X2 \M0/stage1/FA1_0/HA1/_1_  (.A(\M0/prodm1 [0]),
    .B(\M0/prodm2 [0]),
    .Z(\M0/stage1/FA1_0/ha1_sum ));
 AND2_X1 \M0/stage1/FA1_0/HA2/_0_  (.A1(\M0/stage1/FA1_0/ha1_sum ),
    .A2(\M0/stage1/_03_ ),
    .ZN(\M0/stage1/FA1_0/ha2_carry ));
 XOR2_X1 \M0/stage1/FA1_0/HA2/_1_  (.A(\M0/stage1/FA1_0/ha1_sum ),
    .B(\M0/stage1/_03_ ),
    .Z(\M0/stage1/sum1 [0]));
 OR2_X1 \M0/stage1/FA1_0/_0_  (.A1(\M0/stage1/FA1_0/ha1_carry ),
    .A2(\M0/stage1/FA1_0/ha2_carry ),
    .ZN(\M0/stage1/carry1 [0]));
 AND2_X1 \M0/stage1/HA0_0/_0_  (.A1(\M0/prodm1 [0]),
    .A2(\M0/prodm2 [0]),
    .ZN(\M0/stage1/carry0 [0]));
 XOR2_X1 \M0/stage1/HA0_0/_1_  (.A(\M0/prodm1 [0]),
    .B(\M0/prodm2 [0]),
    .Z(\M0/stage1/sum0 [0]));
 INV_X2 \M0/stage1/_04_  (.A(ground),
    .ZN(\M0/stage1/_03_ ));
 MUX2_X2 \M0/stage1/_05_  (.A(\M0/stage1/sum0 [0]),
    .B(\M0/stage1/sum1 [0]),
    .S(ground),
    .Z(\M0/sums1 [0]));
 MUX2_X1 \M0/stage1/_06_  (.A(\M0/stage1/carry0 [0]),
    .B(\M0/stage1/carry1 [0]),
    .S(ground),
    .Z(\M0/stage1/_00_ ));
 MUX2_X2 \M0/stage1/_07_  (.A(\M0/stage1/sum0 [1]),
    .B(\M0/stage1/sum1 [1]),
    .S(\M0/stage1/_00_ ),
    .Z(\M0/sums1 [1]));
 MUX2_X1 \M0/stage1/_08_  (.A(\M0/stage1/carry0 [1]),
    .B(\M0/stage1/carry1 [1]),
    .S(\M0/stage1/_00_ ),
    .Z(\M0/stage1/_01_ ));
 MUX2_X2 \M0/stage1/_09_  (.A(\M0/stage1/sum0 [2]),
    .B(\M0/stage1/sum1 [2]),
    .S(\M0/stage1/_01_ ),
    .Z(\M0/sums1 [2]));
 MUX2_X1 \M0/stage1/_10_  (.A(\M0/stage1/carry0 [2]),
    .B(\M0/stage1/carry1 [2]),
    .S(\M0/stage1/_01_ ),
    .Z(\M0/stage1/_02_ ));
 MUX2_X2 \M0/stage1/_11_  (.A(\M0/stage1/sum0 [3]),
    .B(\M0/stage1/sum1 [3]),
    .S(\M0/stage1/_02_ ),
    .Z(\M0/sums1 [3]));
 MUX2_X1 \M0/stage1/_12_  (.A(\M0/stage1/carry0 [3]),
    .B(\M0/stage1/carry1 [3]),
    .S(\M0/stage1/_02_ ),
    .Z(\M0/c1 ));
 AND2_X1 \M0/stage1/gen_csa[1].FA0/HA1/_0_  (.A1(\M0/prodm1 [1]),
    .A2(\M0/prodm2 [1]),
    .ZN(\M0/stage1/gen_csa[1].FA0/ha1_carry ));
 XOR2_X2 \M0/stage1/gen_csa[1].FA0/HA1/_1_  (.A(\M0/prodm1 [1]),
    .B(\M0/prodm2 [1]),
    .Z(\M0/stage1/gen_csa[1].FA0/ha1_sum ));
 AND2_X1 \M0/stage1/gen_csa[1].FA0/HA2/_0_  (.A1(\M0/stage1/gen_csa[1].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M0/stage1/gen_csa[1].FA0/ha2_carry ));
 XOR2_X1 \M0/stage1/gen_csa[1].FA0/HA2/_1_  (.A(\M0/stage1/gen_csa[1].FA0/ha1_sum ),
    .B(ground),
    .Z(\M0/stage1/sum0 [1]));
 OR2_X1 \M0/stage1/gen_csa[1].FA0/_0_  (.A1(\M0/stage1/gen_csa[1].FA0/ha1_carry ),
    .A2(\M0/stage1/gen_csa[1].FA0/ha2_carry ),
    .ZN(\M0/stage1/carry0 [1]));
 AND2_X1 \M0/stage1/gen_csa[1].FA1/HA1/_0_  (.A1(\M0/prodm1 [1]),
    .A2(\M0/prodm2 [1]),
    .ZN(\M0/stage1/gen_csa[1].FA1/ha1_carry ));
 XOR2_X2 \M0/stage1/gen_csa[1].FA1/HA1/_1_  (.A(\M0/prodm1 [1]),
    .B(\M0/prodm2 [1]),
    .Z(\M0/stage1/gen_csa[1].FA1/ha1_sum ));
 AND2_X1 \M0/stage1/gen_csa[1].FA1/HA2/_0_  (.A1(\M0/stage1/gen_csa[1].FA1/ha1_sum ),
    .A2(\M0/stage1/_03_ ),
    .ZN(\M0/stage1/gen_csa[1].FA1/ha2_carry ));
 XOR2_X1 \M0/stage1/gen_csa[1].FA1/HA2/_1_  (.A(\M0/stage1/gen_csa[1].FA1/ha1_sum ),
    .B(\M0/stage1/_03_ ),
    .Z(\M0/stage1/sum1 [1]));
 OR2_X1 \M0/stage1/gen_csa[1].FA1/_0_  (.A1(\M0/stage1/gen_csa[1].FA1/ha1_carry ),
    .A2(\M0/stage1/gen_csa[1].FA1/ha2_carry ),
    .ZN(\M0/stage1/carry1 [1]));
 AND2_X1 \M0/stage1/gen_csa[2].FA0/HA1/_0_  (.A1(\M0/prodm1 [2]),
    .A2(\M0/prodm2 [2]),
    .ZN(\M0/stage1/gen_csa[2].FA0/ha1_carry ));
 XOR2_X2 \M0/stage1/gen_csa[2].FA0/HA1/_1_  (.A(\M0/prodm1 [2]),
    .B(\M0/prodm2 [2]),
    .Z(\M0/stage1/gen_csa[2].FA0/ha1_sum ));
 AND2_X1 \M0/stage1/gen_csa[2].FA0/HA2/_0_  (.A1(\M0/stage1/gen_csa[2].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M0/stage1/gen_csa[2].FA0/ha2_carry ));
 XOR2_X1 \M0/stage1/gen_csa[2].FA0/HA2/_1_  (.A(\M0/stage1/gen_csa[2].FA0/ha1_sum ),
    .B(ground),
    .Z(\M0/stage1/sum0 [2]));
 OR2_X1 \M0/stage1/gen_csa[2].FA0/_0_  (.A1(\M0/stage1/gen_csa[2].FA0/ha1_carry ),
    .A2(\M0/stage1/gen_csa[2].FA0/ha2_carry ),
    .ZN(\M0/stage1/carry0 [2]));
 AND2_X1 \M0/stage1/gen_csa[2].FA1/HA1/_0_  (.A1(\M0/prodm1 [2]),
    .A2(\M0/prodm2 [2]),
    .ZN(\M0/stage1/gen_csa[2].FA1/ha1_carry ));
 XOR2_X2 \M0/stage1/gen_csa[2].FA1/HA1/_1_  (.A(\M0/prodm1 [2]),
    .B(\M0/prodm2 [2]),
    .Z(\M0/stage1/gen_csa[2].FA1/ha1_sum ));
 AND2_X1 \M0/stage1/gen_csa[2].FA1/HA2/_0_  (.A1(\M0/stage1/gen_csa[2].FA1/ha1_sum ),
    .A2(\M0/stage1/_03_ ),
    .ZN(\M0/stage1/gen_csa[2].FA1/ha2_carry ));
 XOR2_X1 \M0/stage1/gen_csa[2].FA1/HA2/_1_  (.A(\M0/stage1/gen_csa[2].FA1/ha1_sum ),
    .B(\M0/stage1/_03_ ),
    .Z(\M0/stage1/sum1 [2]));
 OR2_X1 \M0/stage1/gen_csa[2].FA1/_0_  (.A1(\M0/stage1/gen_csa[2].FA1/ha1_carry ),
    .A2(\M0/stage1/gen_csa[2].FA1/ha2_carry ),
    .ZN(\M0/stage1/carry1 [2]));
 AND2_X1 \M0/stage1/gen_csa[3].FA0/HA1/_0_  (.A1(\M0/prodm1 [3]),
    .A2(\M0/prodm2 [3]),
    .ZN(\M0/stage1/gen_csa[3].FA0/ha1_carry ));
 XOR2_X2 \M0/stage1/gen_csa[3].FA0/HA1/_1_  (.A(\M0/prodm1 [3]),
    .B(\M0/prodm2 [3]),
    .Z(\M0/stage1/gen_csa[3].FA0/ha1_sum ));
 AND2_X1 \M0/stage1/gen_csa[3].FA0/HA2/_0_  (.A1(\M0/stage1/gen_csa[3].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M0/stage1/gen_csa[3].FA0/ha2_carry ));
 XOR2_X1 \M0/stage1/gen_csa[3].FA0/HA2/_1_  (.A(\M0/stage1/gen_csa[3].FA0/ha1_sum ),
    .B(ground),
    .Z(\M0/stage1/sum0 [3]));
 OR2_X1 \M0/stage1/gen_csa[3].FA0/_0_  (.A1(\M0/stage1/gen_csa[3].FA0/ha1_carry ),
    .A2(\M0/stage1/gen_csa[3].FA0/ha2_carry ),
    .ZN(\M0/stage1/carry0 [3]));
 AND2_X1 \M0/stage1/gen_csa[3].FA1/HA1/_0_  (.A1(\M0/prodm1 [3]),
    .A2(\M0/prodm2 [3]),
    .ZN(\M0/stage1/gen_csa[3].FA1/ha1_carry ));
 XOR2_X2 \M0/stage1/gen_csa[3].FA1/HA1/_1_  (.A(\M0/prodm1 [3]),
    .B(\M0/prodm2 [3]),
    .Z(\M0/stage1/gen_csa[3].FA1/ha1_sum ));
 AND2_X1 \M0/stage1/gen_csa[3].FA1/HA2/_0_  (.A1(\M0/stage1/gen_csa[3].FA1/ha1_sum ),
    .A2(\M0/stage1/_03_ ),
    .ZN(\M0/stage1/gen_csa[3].FA1/ha2_carry ));
 XOR2_X1 \M0/stage1/gen_csa[3].FA1/HA2/_1_  (.A(\M0/stage1/gen_csa[3].FA1/ha1_sum ),
    .B(\M0/stage1/_03_ ),
    .Z(\M0/stage1/sum1 [3]));
 OR2_X1 \M0/stage1/gen_csa[3].FA1/_0_  (.A1(\M0/stage1/gen_csa[3].FA1/ha1_carry ),
    .A2(\M0/stage1/gen_csa[3].FA1/ha2_carry ),
    .ZN(\M0/stage1/carry1 [3]));
 AND2_X1 \M0/stage2/FA1_0/HA1/_0_  (.A1(\M0/prodm0 [2]),
    .A2(\M0/sums1 [0]),
    .ZN(\M0/stage2/FA1_0/ha1_carry ));
 XOR2_X2 \M0/stage2/FA1_0/HA1/_1_  (.A(\M0/prodm0 [2]),
    .B(\M0/sums1 [0]),
    .Z(\M0/stage2/FA1_0/ha1_sum ));
 AND2_X1 \M0/stage2/FA1_0/HA2/_0_  (.A1(\M0/stage2/FA1_0/ha1_sum ),
    .A2(\M0/stage2/_03_ ),
    .ZN(\M0/stage2/FA1_0/ha2_carry ));
 XOR2_X1 \M0/stage2/FA1_0/HA2/_1_  (.A(\M0/stage2/FA1_0/ha1_sum ),
    .B(\M0/stage2/_03_ ),
    .Z(\M0/stage2/sum1 [0]));
 OR2_X1 \M0/stage2/FA1_0/_0_  (.A1(\M0/stage2/FA1_0/ha1_carry ),
    .A2(\M0/stage2/FA1_0/ha2_carry ),
    .ZN(\M0/stage2/carry1 [0]));
 AND2_X1 \M0/stage2/HA0_0/_0_  (.A1(\M0/prodm0 [2]),
    .A2(\M0/sums1 [0]),
    .ZN(\M0/stage2/carry0 [0]));
 XOR2_X1 \M0/stage2/HA0_0/_1_  (.A(\M0/prodm0 [2]),
    .B(\M0/sums1 [0]),
    .Z(\M0/stage2/sum0 [0]));
 INV_X2 \M0/stage2/_04_  (.A(ground),
    .ZN(\M0/stage2/_03_ ));
 MUX2_X1 \M0/stage2/_05_  (.A(\M0/stage2/sum0 [0]),
    .B(\M0/stage2/sum1 [0]),
    .S(ground),
    .Z(prodm0[2]));
 MUX2_X1 \M0/stage2/_06_  (.A(\M0/stage2/carry0 [0]),
    .B(\M0/stage2/carry1 [0]),
    .S(ground),
    .Z(\M0/stage2/_00_ ));
 MUX2_X1 \M0/stage2/_07_  (.A(\M0/stage2/sum0 [1]),
    .B(\M0/stage2/sum1 [1]),
    .S(\M0/stage2/_00_ ),
    .Z(prodm0[3]));
 MUX2_X1 \M0/stage2/_08_  (.A(\M0/stage2/carry0 [1]),
    .B(\M0/stage2/carry1 [1]),
    .S(\M0/stage2/_00_ ),
    .Z(\M0/stage2/_01_ ));
 MUX2_X2 \M0/stage2/_09_  (.A(\M0/stage2/sum0 [2]),
    .B(\M0/stage2/sum1 [2]),
    .S(\M0/stage2/_01_ ),
    .Z(\M0/sums2 [2]));
 MUX2_X1 \M0/stage2/_10_  (.A(\M0/stage2/carry0 [2]),
    .B(\M0/stage2/carry1 [2]),
    .S(\M0/stage2/_01_ ),
    .Z(\M0/stage2/_02_ ));
 MUX2_X2 \M0/stage2/_11_  (.A(\M0/stage2/sum0 [3]),
    .B(\M0/stage2/sum1 [3]),
    .S(\M0/stage2/_02_ ),
    .Z(\M0/sums2 [3]));
 MUX2_X1 \M0/stage2/_12_  (.A(\M0/stage2/carry0 [3]),
    .B(\M0/stage2/carry1 [3]),
    .S(\M0/stage2/_02_ ),
    .Z(\M0/c2 ));
 AND2_X1 \M0/stage2/gen_csa[1].FA0/HA1/_0_  (.A1(\M0/prodm0 [3]),
    .A2(\M0/sums1 [1]),
    .ZN(\M0/stage2/gen_csa[1].FA0/ha1_carry ));
 XOR2_X2 \M0/stage2/gen_csa[1].FA0/HA1/_1_  (.A(\M0/prodm0 [3]),
    .B(\M0/sums1 [1]),
    .Z(\M0/stage2/gen_csa[1].FA0/ha1_sum ));
 AND2_X1 \M0/stage2/gen_csa[1].FA0/HA2/_0_  (.A1(\M0/stage2/gen_csa[1].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M0/stage2/gen_csa[1].FA0/ha2_carry ));
 XOR2_X1 \M0/stage2/gen_csa[1].FA0/HA2/_1_  (.A(\M0/stage2/gen_csa[1].FA0/ha1_sum ),
    .B(ground),
    .Z(\M0/stage2/sum0 [1]));
 OR2_X1 \M0/stage2/gen_csa[1].FA0/_0_  (.A1(\M0/stage2/gen_csa[1].FA0/ha1_carry ),
    .A2(\M0/stage2/gen_csa[1].FA0/ha2_carry ),
    .ZN(\M0/stage2/carry0 [1]));
 AND2_X1 \M0/stage2/gen_csa[1].FA1/HA1/_0_  (.A1(\M0/prodm0 [3]),
    .A2(\M0/sums1 [1]),
    .ZN(\M0/stage2/gen_csa[1].FA1/ha1_carry ));
 XOR2_X2 \M0/stage2/gen_csa[1].FA1/HA1/_1_  (.A(\M0/prodm0 [3]),
    .B(\M0/sums1 [1]),
    .Z(\M0/stage2/gen_csa[1].FA1/ha1_sum ));
 AND2_X1 \M0/stage2/gen_csa[1].FA1/HA2/_0_  (.A1(\M0/stage2/gen_csa[1].FA1/ha1_sum ),
    .A2(\M0/stage2/_03_ ),
    .ZN(\M0/stage2/gen_csa[1].FA1/ha2_carry ));
 XOR2_X1 \M0/stage2/gen_csa[1].FA1/HA2/_1_  (.A(\M0/stage2/gen_csa[1].FA1/ha1_sum ),
    .B(\M0/stage2/_03_ ),
    .Z(\M0/stage2/sum1 [1]));
 OR2_X1 \M0/stage2/gen_csa[1].FA1/_0_  (.A1(\M0/stage2/gen_csa[1].FA1/ha1_carry ),
    .A2(\M0/stage2/gen_csa[1].FA1/ha2_carry ),
    .ZN(\M0/stage2/carry1 [1]));
 AND2_X1 \M0/stage2/gen_csa[2].FA0/HA1/_0_  (.A1(ground),
    .A2(\M0/sums1 [2]),
    .ZN(\M0/stage2/gen_csa[2].FA0/ha1_carry ));
 XOR2_X2 \M0/stage2/gen_csa[2].FA0/HA1/_1_  (.A(ground),
    .B(\M0/sums1 [2]),
    .Z(\M0/stage2/gen_csa[2].FA0/ha1_sum ));
 AND2_X1 \M0/stage2/gen_csa[2].FA0/HA2/_0_  (.A1(\M0/stage2/gen_csa[2].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M0/stage2/gen_csa[2].FA0/ha2_carry ));
 XOR2_X1 \M0/stage2/gen_csa[2].FA0/HA2/_1_  (.A(\M0/stage2/gen_csa[2].FA0/ha1_sum ),
    .B(ground),
    .Z(\M0/stage2/sum0 [2]));
 OR2_X1 \M0/stage2/gen_csa[2].FA0/_0_  (.A1(\M0/stage2/gen_csa[2].FA0/ha1_carry ),
    .A2(\M0/stage2/gen_csa[2].FA0/ha2_carry ),
    .ZN(\M0/stage2/carry0 [2]));
 AND2_X1 \M0/stage2/gen_csa[2].FA1/HA1/_0_  (.A1(ground),
    .A2(\M0/sums1 [2]),
    .ZN(\M0/stage2/gen_csa[2].FA1/ha1_carry ));
 XOR2_X2 \M0/stage2/gen_csa[2].FA1/HA1/_1_  (.A(ground),
    .B(\M0/sums1 [2]),
    .Z(\M0/stage2/gen_csa[2].FA1/ha1_sum ));
 AND2_X1 \M0/stage2/gen_csa[2].FA1/HA2/_0_  (.A1(\M0/stage2/gen_csa[2].FA1/ha1_sum ),
    .A2(\M0/stage2/_03_ ),
    .ZN(\M0/stage2/gen_csa[2].FA1/ha2_carry ));
 XOR2_X1 \M0/stage2/gen_csa[2].FA1/HA2/_1_  (.A(\M0/stage2/gen_csa[2].FA1/ha1_sum ),
    .B(\M0/stage2/_03_ ),
    .Z(\M0/stage2/sum1 [2]));
 OR2_X1 \M0/stage2/gen_csa[2].FA1/_0_  (.A1(\M0/stage2/gen_csa[2].FA1/ha1_carry ),
    .A2(\M0/stage2/gen_csa[2].FA1/ha2_carry ),
    .ZN(\M0/stage2/carry1 [2]));
 AND2_X1 \M0/stage2/gen_csa[3].FA0/HA1/_0_  (.A1(ground),
    .A2(\M0/sums1 [3]),
    .ZN(\M0/stage2/gen_csa[3].FA0/ha1_carry ));
 XOR2_X2 \M0/stage2/gen_csa[3].FA0/HA1/_1_  (.A(ground),
    .B(\M0/sums1 [3]),
    .Z(\M0/stage2/gen_csa[3].FA0/ha1_sum ));
 AND2_X1 \M0/stage2/gen_csa[3].FA0/HA2/_0_  (.A1(\M0/stage2/gen_csa[3].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M0/stage2/gen_csa[3].FA0/ha2_carry ));
 XOR2_X1 \M0/stage2/gen_csa[3].FA0/HA2/_1_  (.A(\M0/stage2/gen_csa[3].FA0/ha1_sum ),
    .B(ground),
    .Z(\M0/stage2/sum0 [3]));
 OR2_X1 \M0/stage2/gen_csa[3].FA0/_0_  (.A1(\M0/stage2/gen_csa[3].FA0/ha1_carry ),
    .A2(\M0/stage2/gen_csa[3].FA0/ha2_carry ),
    .ZN(\M0/stage2/carry0 [3]));
 AND2_X1 \M0/stage2/gen_csa[3].FA1/HA1/_0_  (.A1(ground),
    .A2(\M0/sums1 [3]),
    .ZN(\M0/stage2/gen_csa[3].FA1/ha1_carry ));
 XOR2_X2 \M0/stage2/gen_csa[3].FA1/HA1/_1_  (.A(ground),
    .B(\M0/sums1 [3]),
    .Z(\M0/stage2/gen_csa[3].FA1/ha1_sum ));
 AND2_X1 \M0/stage2/gen_csa[3].FA1/HA2/_0_  (.A1(\M0/stage2/gen_csa[3].FA1/ha1_sum ),
    .A2(\M0/stage2/_03_ ),
    .ZN(\M0/stage2/gen_csa[3].FA1/ha2_carry ));
 XOR2_X1 \M0/stage2/gen_csa[3].FA1/HA2/_1_  (.A(\M0/stage2/gen_csa[3].FA1/ha1_sum ),
    .B(\M0/stage2/_03_ ),
    .Z(\M0/stage2/sum1 [3]));
 OR2_X1 \M0/stage2/gen_csa[3].FA1/_0_  (.A1(\M0/stage2/gen_csa[3].FA1/ha1_carry ),
    .A2(\M0/stage2/gen_csa[3].FA1/ha2_carry ),
    .ZN(\M0/stage2/carry1 [3]));
 AND2_X1 \M0/stage3/FA1_0/HA1/_0_  (.A1(\M0/sums2 [2]),
    .A2(\M0/prodm3 [0]),
    .ZN(\M0/stage3/FA1_0/ha1_carry ));
 XOR2_X2 \M0/stage3/FA1_0/HA1/_1_  (.A(\M0/sums2 [2]),
    .B(\M0/prodm3 [0]),
    .Z(\M0/stage3/FA1_0/ha1_sum ));
 AND2_X1 \M0/stage3/FA1_0/HA2/_0_  (.A1(\M0/stage3/FA1_0/ha1_sum ),
    .A2(\M0/stage3/_03_ ),
    .ZN(\M0/stage3/FA1_0/ha2_carry ));
 XOR2_X1 \M0/stage3/FA1_0/HA2/_1_  (.A(\M0/stage3/FA1_0/ha1_sum ),
    .B(\M0/stage3/_03_ ),
    .Z(\M0/stage3/sum1 [0]));
 OR2_X1 \M0/stage3/FA1_0/_0_  (.A1(\M0/stage3/FA1_0/ha1_carry ),
    .A2(\M0/stage3/FA1_0/ha2_carry ),
    .ZN(\M0/stage3/carry1 [0]));
 AND2_X1 \M0/stage3/HA0_0/_0_  (.A1(\M0/sums2 [2]),
    .A2(\M0/prodm3 [0]),
    .ZN(\M0/stage3/carry0 [0]));
 XOR2_X1 \M0/stage3/HA0_0/_1_  (.A(\M0/sums2 [2]),
    .B(\M0/prodm3 [0]),
    .Z(\M0/stage3/sum0 [0]));
 INV_X2 \M0/stage3/_04_  (.A(ground),
    .ZN(\M0/stage3/_03_ ));
 MUX2_X1 \M0/stage3/_05_  (.A(\M0/stage3/sum0 [0]),
    .B(\M0/stage3/sum1 [0]),
    .S(ground),
    .Z(prodm0[4]));
 MUX2_X1 \M0/stage3/_06_  (.A(\M0/stage3/carry0 [0]),
    .B(\M0/stage3/carry1 [0]),
    .S(ground),
    .Z(\M0/stage3/_00_ ));
 MUX2_X1 \M0/stage3/_07_  (.A(\M0/stage3/sum0 [1]),
    .B(\M0/stage3/sum1 [1]),
    .S(\M0/stage3/_00_ ),
    .Z(prodm0[5]));
 MUX2_X1 \M0/stage3/_08_  (.A(\M0/stage3/carry0 [1]),
    .B(\M0/stage3/carry1 [1]),
    .S(\M0/stage3/_00_ ),
    .Z(\M0/stage3/_01_ ));
 MUX2_X1 \M0/stage3/_09_  (.A(\M0/stage3/sum0 [2]),
    .B(\M0/stage3/sum1 [2]),
    .S(\M0/stage3/_01_ ),
    .Z(prodm0[6]));
 MUX2_X1 \M0/stage3/_10_  (.A(\M0/stage3/carry0 [2]),
    .B(\M0/stage3/carry1 [2]),
    .S(\M0/stage3/_01_ ),
    .Z(\M0/stage3/_02_ ));
 MUX2_X1 \M0/stage3/_11_  (.A(\M0/stage3/sum0 [3]),
    .B(\M0/stage3/sum1 [3]),
    .S(\M0/stage3/_02_ ),
    .Z(prodm0[7]));
 MUX2_X1 \M0/stage3/_12_  (.A(\M0/stage3/carry0 [3]),
    .B(\M0/stage3/carry1 [3]),
    .S(\M0/stage3/_02_ ),
    .Z(ov1));
 AND2_X1 \M0/stage3/gen_csa[1].FA0/HA1/_0_  (.A1(\M0/sums2 [3]),
    .A2(\M0/prodm3 [1]),
    .ZN(\M0/stage3/gen_csa[1].FA0/ha1_carry ));
 XOR2_X2 \M0/stage3/gen_csa[1].FA0/HA1/_1_  (.A(\M0/sums2 [3]),
    .B(\M0/prodm3 [1]),
    .Z(\M0/stage3/gen_csa[1].FA0/ha1_sum ));
 AND2_X1 \M0/stage3/gen_csa[1].FA0/HA2/_0_  (.A1(\M0/stage3/gen_csa[1].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M0/stage3/gen_csa[1].FA0/ha2_carry ));
 XOR2_X1 \M0/stage3/gen_csa[1].FA0/HA2/_1_  (.A(\M0/stage3/gen_csa[1].FA0/ha1_sum ),
    .B(ground),
    .Z(\M0/stage3/sum0 [1]));
 OR2_X1 \M0/stage3/gen_csa[1].FA0/_0_  (.A1(\M0/stage3/gen_csa[1].FA0/ha1_carry ),
    .A2(\M0/stage3/gen_csa[1].FA0/ha2_carry ),
    .ZN(\M0/stage3/carry0 [1]));
 AND2_X1 \M0/stage3/gen_csa[1].FA1/HA1/_0_  (.A1(\M0/sums2 [3]),
    .A2(\M0/prodm3 [1]),
    .ZN(\M0/stage3/gen_csa[1].FA1/ha1_carry ));
 XOR2_X2 \M0/stage3/gen_csa[1].FA1/HA1/_1_  (.A(\M0/sums2 [3]),
    .B(\M0/prodm3 [1]),
    .Z(\M0/stage3/gen_csa[1].FA1/ha1_sum ));
 AND2_X1 \M0/stage3/gen_csa[1].FA1/HA2/_0_  (.A1(\M0/stage3/gen_csa[1].FA1/ha1_sum ),
    .A2(\M0/stage3/_03_ ),
    .ZN(\M0/stage3/gen_csa[1].FA1/ha2_carry ));
 XOR2_X1 \M0/stage3/gen_csa[1].FA1/HA2/_1_  (.A(\M0/stage3/gen_csa[1].FA1/ha1_sum ),
    .B(\M0/stage3/_03_ ),
    .Z(\M0/stage3/sum1 [1]));
 OR2_X1 \M0/stage3/gen_csa[1].FA1/_0_  (.A1(\M0/stage3/gen_csa[1].FA1/ha1_carry ),
    .A2(\M0/stage3/gen_csa[1].FA1/ha2_carry ),
    .ZN(\M0/stage3/carry1 [1]));
 AND2_X1 \M0/stage3/gen_csa[2].FA0/HA1/_0_  (.A1(\M0/cnet ),
    .A2(\M0/prodm3 [2]),
    .ZN(\M0/stage3/gen_csa[2].FA0/ha1_carry ));
 XOR2_X2 \M0/stage3/gen_csa[2].FA0/HA1/_1_  (.A(\M0/cnet ),
    .B(\M0/prodm3 [2]),
    .Z(\M0/stage3/gen_csa[2].FA0/ha1_sum ));
 AND2_X1 \M0/stage3/gen_csa[2].FA0/HA2/_0_  (.A1(\M0/stage3/gen_csa[2].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M0/stage3/gen_csa[2].FA0/ha2_carry ));
 XOR2_X1 \M0/stage3/gen_csa[2].FA0/HA2/_1_  (.A(\M0/stage3/gen_csa[2].FA0/ha1_sum ),
    .B(ground),
    .Z(\M0/stage3/sum0 [2]));
 OR2_X1 \M0/stage3/gen_csa[2].FA0/_0_  (.A1(\M0/stage3/gen_csa[2].FA0/ha1_carry ),
    .A2(\M0/stage3/gen_csa[2].FA0/ha2_carry ),
    .ZN(\M0/stage3/carry0 [2]));
 AND2_X1 \M0/stage3/gen_csa[2].FA1/HA1/_0_  (.A1(\M0/cnet ),
    .A2(\M0/prodm3 [2]),
    .ZN(\M0/stage3/gen_csa[2].FA1/ha1_carry ));
 XOR2_X2 \M0/stage3/gen_csa[2].FA1/HA1/_1_  (.A(\M0/cnet ),
    .B(\M0/prodm3 [2]),
    .Z(\M0/stage3/gen_csa[2].FA1/ha1_sum ));
 AND2_X1 \M0/stage3/gen_csa[2].FA1/HA2/_0_  (.A1(\M0/stage3/gen_csa[2].FA1/ha1_sum ),
    .A2(\M0/stage3/_03_ ),
    .ZN(\M0/stage3/gen_csa[2].FA1/ha2_carry ));
 XOR2_X1 \M0/stage3/gen_csa[2].FA1/HA2/_1_  (.A(\M0/stage3/gen_csa[2].FA1/ha1_sum ),
    .B(\M0/stage3/_03_ ),
    .Z(\M0/stage3/sum1 [2]));
 OR2_X1 \M0/stage3/gen_csa[2].FA1/_0_  (.A1(\M0/stage3/gen_csa[2].FA1/ha1_carry ),
    .A2(\M0/stage3/gen_csa[2].FA1/ha2_carry ),
    .ZN(\M0/stage3/carry1 [2]));
 AND2_X1 \M0/stage3/gen_csa[3].FA0/HA1/_0_  (.A1(ground),
    .A2(\M0/prodm3 [3]),
    .ZN(\M0/stage3/gen_csa[3].FA0/ha1_carry ));
 XOR2_X2 \M0/stage3/gen_csa[3].FA0/HA1/_1_  (.A(ground),
    .B(\M0/prodm3 [3]),
    .Z(\M0/stage3/gen_csa[3].FA0/ha1_sum ));
 AND2_X1 \M0/stage3/gen_csa[3].FA0/HA2/_0_  (.A1(\M0/stage3/gen_csa[3].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M0/stage3/gen_csa[3].FA0/ha2_carry ));
 XOR2_X1 \M0/stage3/gen_csa[3].FA0/HA2/_1_  (.A(\M0/stage3/gen_csa[3].FA0/ha1_sum ),
    .B(ground),
    .Z(\M0/stage3/sum0 [3]));
 OR2_X1 \M0/stage3/gen_csa[3].FA0/_0_  (.A1(\M0/stage3/gen_csa[3].FA0/ha1_carry ),
    .A2(\M0/stage3/gen_csa[3].FA0/ha2_carry ),
    .ZN(\M0/stage3/carry0 [3]));
 AND2_X1 \M0/stage3/gen_csa[3].FA1/HA1/_0_  (.A1(ground),
    .A2(\M0/prodm3 [3]),
    .ZN(\M0/stage3/gen_csa[3].FA1/ha1_carry ));
 XOR2_X1 \M0/stage3/gen_csa[3].FA1/HA1/_1_  (.A(ground),
    .B(\M0/prodm3 [3]),
    .Z(\M0/stage3/gen_csa[3].FA1/ha1_sum ));
 AND2_X1 \M0/stage3/gen_csa[3].FA1/HA2/_0_  (.A1(\M0/stage3/gen_csa[3].FA1/ha1_sum ),
    .A2(\M0/stage3/_03_ ),
    .ZN(\M0/stage3/gen_csa[3].FA1/ha2_carry ));
 XOR2_X1 \M0/stage3/gen_csa[3].FA1/HA2/_1_  (.A(\M0/stage3/gen_csa[3].FA1/ha1_sum ),
    .B(\M0/stage3/_03_ ),
    .Z(\M0/stage3/sum1 [3]));
 OR2_X1 \M0/stage3/gen_csa[3].FA1/_0_  (.A1(\M0/stage3/gen_csa[3].FA1/ha1_carry ),
    .A2(\M0/stage3/gen_csa[3].FA1/ha2_carry ),
    .ZN(\M0/stage3/carry1 [3]));
 AND2_X1 \M1/M0/HA0/_0_  (.A1(\M1/M0/a0b1 ),
    .A2(\M1/M0/a1b0 ),
    .ZN(\M1/M0/carry ));
 XOR2_X1 \M1/M0/HA0/_1_  (.A(\M1/M0/a0b1 ),
    .B(\M1/M0/a1b0 ),
    .Z(prodm1[1]));
 AND2_X1 \M1/M0/HA1/_0_  (.A1(\M1/M0/a1b1 ),
    .A2(\M1/M0/carry ),
    .ZN(\M1/prodm0 [3]));
 XOR2_X2 \M1/M0/HA1/_1_  (.A(\M1/M0/a1b1 ),
    .B(\M1/M0/carry ),
    .Z(\M1/prodm0 [2]));
 AND2_X1 \M1/M0/_0_  (.A1(a[1]),
    .A2(b[5]),
    .ZN(\M1/M0/a1b1 ));
 AND2_X1 \M1/M0/_1_  (.A1(b[5]),
    .A2(a[0]),
    .ZN(\M1/M0/a0b1 ));
 AND2_X1 \M1/M0/_2_  (.A1(a[1]),
    .A2(b[4]),
    .ZN(\M1/M0/a1b0 ));
 AND2_X1 \M1/M0/_3_  (.A1(a[0]),
    .A2(b[4]),
    .ZN(prodm1[0]));
 AND2_X1 \M1/M1/HA0/_0_  (.A1(\M1/M1/a0b1 ),
    .A2(\M1/M1/a1b0 ),
    .ZN(\M1/M1/carry ));
 XOR2_X2 \M1/M1/HA0/_1_  (.A(\M1/M1/a0b1 ),
    .B(\M1/M1/a1b0 ),
    .Z(\M1/prodm1 [1]));
 AND2_X2 \M1/M1/HA1/_0_  (.A1(\M1/M1/a1b1 ),
    .A2(\M1/M1/carry ),
    .ZN(\M1/prodm1 [3]));
 XOR2_X2 \M1/M1/HA1/_1_  (.A(\M1/M1/a1b1 ),
    .B(\M1/M1/carry ),
    .Z(\M1/prodm1 [2]));
 AND2_X1 \M1/M1/_0_  (.A1(a[1]),
    .A2(b[7]),
    .ZN(\M1/M1/a1b1 ));
 AND2_X1 \M1/M1/_1_  (.A1(b[7]),
    .A2(a[0]),
    .ZN(\M1/M1/a0b1 ));
 AND2_X1 \M1/M1/_2_  (.A1(a[1]),
    .A2(b[6]),
    .ZN(\M1/M1/a1b0 ));
 AND2_X1 \M1/M1/_3_  (.A1(a[0]),
    .A2(b[6]),
    .ZN(\M1/prodm1 [0]));
 AND2_X1 \M1/M2/HA0/_0_  (.A1(\M1/M2/a0b1 ),
    .A2(\M1/M2/a1b0 ),
    .ZN(\M1/M2/carry ));
 XOR2_X2 \M1/M2/HA0/_1_  (.A(\M1/M2/a0b1 ),
    .B(\M1/M2/a1b0 ),
    .Z(\M1/prodm2 [1]));
 AND2_X2 \M1/M2/HA1/_0_  (.A1(\M1/M2/a1b1 ),
    .A2(\M1/M2/carry ),
    .ZN(\M1/prodm2 [3]));
 XOR2_X2 \M1/M2/HA1/_1_  (.A(\M1/M2/a1b1 ),
    .B(\M1/M2/carry ),
    .Z(\M1/prodm2 [2]));
 AND2_X1 \M1/M2/_0_  (.A1(a[3]),
    .A2(b[5]),
    .ZN(\M1/M2/a1b1 ));
 AND2_X1 \M1/M2/_1_  (.A1(b[5]),
    .A2(a[2]),
    .ZN(\M1/M2/a0b1 ));
 AND2_X1 \M1/M2/_2_  (.A1(a[3]),
    .A2(b[4]),
    .ZN(\M1/M2/a1b0 ));
 AND2_X1 \M1/M2/_3_  (.A1(a[2]),
    .A2(b[4]),
    .ZN(\M1/prodm2 [0]));
 AND2_X1 \M1/M3/HA0/_0_  (.A1(\M1/M3/a0b1 ),
    .A2(\M1/M3/a1b0 ),
    .ZN(\M1/M3/carry ));
 XOR2_X2 \M1/M3/HA0/_1_  (.A(\M1/M3/a0b1 ),
    .B(\M1/M3/a1b0 ),
    .Z(\M1/prodm3 [1]));
 AND2_X1 \M1/M3/HA1/_0_  (.A1(\M1/M3/a1b1 ),
    .A2(\M1/M3/carry ),
    .ZN(\M1/prodm3 [3]));
 XOR2_X2 \M1/M3/HA1/_1_  (.A(\M1/M3/a1b1 ),
    .B(\M1/M3/carry ),
    .Z(\M1/prodm3 [2]));
 AND2_X1 \M1/M3/_0_  (.A1(a[3]),
    .A2(b[7]),
    .ZN(\M1/M3/a1b1 ));
 AND2_X1 \M1/M3/_1_  (.A1(b[7]),
    .A2(a[2]),
    .ZN(\M1/M3/a0b1 ));
 AND2_X1 \M1/M3/_2_  (.A1(a[3]),
    .A2(b[6]),
    .ZN(\M1/M3/a1b0 ));
 AND2_X1 \M1/M3/_3_  (.A1(a[2]),
    .A2(b[6]),
    .ZN(\M1/prodm3 [0]));
 OR2_X2 \M1/_0_  (.A1(\M1/c1 ),
    .A2(\M1/c2 ),
    .ZN(\M1/cnet ));
 AND2_X1 \M1/stage1/FA1_0/HA1/_0_  (.A1(\M1/prodm1 [0]),
    .A2(\M1/prodm2 [0]),
    .ZN(\M1/stage1/FA1_0/ha1_carry ));
 XOR2_X2 \M1/stage1/FA1_0/HA1/_1_  (.A(\M1/prodm1 [0]),
    .B(\M1/prodm2 [0]),
    .Z(\M1/stage1/FA1_0/ha1_sum ));
 AND2_X1 \M1/stage1/FA1_0/HA2/_0_  (.A1(\M1/stage1/FA1_0/ha1_sum ),
    .A2(\M1/stage1/_03_ ),
    .ZN(\M1/stage1/FA1_0/ha2_carry ));
 XOR2_X1 \M1/stage1/FA1_0/HA2/_1_  (.A(\M1/stage1/FA1_0/ha1_sum ),
    .B(\M1/stage1/_03_ ),
    .Z(\M1/stage1/sum1 [0]));
 OR2_X1 \M1/stage1/FA1_0/_0_  (.A1(\M1/stage1/FA1_0/ha1_carry ),
    .A2(\M1/stage1/FA1_0/ha2_carry ),
    .ZN(\M1/stage1/carry1 [0]));
 AND2_X1 \M1/stage1/HA0_0/_0_  (.A1(\M1/prodm1 [0]),
    .A2(\M1/prodm2 [0]),
    .ZN(\M1/stage1/carry0 [0]));
 XOR2_X1 \M1/stage1/HA0_0/_1_  (.A(\M1/prodm1 [0]),
    .B(\M1/prodm2 [0]),
    .Z(\M1/stage1/sum0 [0]));
 INV_X2 \M1/stage1/_04_  (.A(ground),
    .ZN(\M1/stage1/_03_ ));
 MUX2_X2 \M1/stage1/_05_  (.A(\M1/stage1/sum0 [0]),
    .B(\M1/stage1/sum1 [0]),
    .S(ground),
    .Z(\M1/sums1 [0]));
 MUX2_X1 \M1/stage1/_06_  (.A(\M1/stage1/carry0 [0]),
    .B(\M1/stage1/carry1 [0]),
    .S(ground),
    .Z(\M1/stage1/_00_ ));
 MUX2_X2 \M1/stage1/_07_  (.A(\M1/stage1/sum0 [1]),
    .B(\M1/stage1/sum1 [1]),
    .S(\M1/stage1/_00_ ),
    .Z(\M1/sums1 [1]));
 MUX2_X1 \M1/stage1/_08_  (.A(\M1/stage1/carry0 [1]),
    .B(\M1/stage1/carry1 [1]),
    .S(\M1/stage1/_00_ ),
    .Z(\M1/stage1/_01_ ));
 MUX2_X2 \M1/stage1/_09_  (.A(\M1/stage1/sum0 [2]),
    .B(\M1/stage1/sum1 [2]),
    .S(\M1/stage1/_01_ ),
    .Z(\M1/sums1 [2]));
 MUX2_X1 \M1/stage1/_10_  (.A(\M1/stage1/carry0 [2]),
    .B(\M1/stage1/carry1 [2]),
    .S(\M1/stage1/_01_ ),
    .Z(\M1/stage1/_02_ ));
 MUX2_X2 \M1/stage1/_11_  (.A(\M1/stage1/sum0 [3]),
    .B(\M1/stage1/sum1 [3]),
    .S(\M1/stage1/_02_ ),
    .Z(\M1/sums1 [3]));
 MUX2_X1 \M1/stage1/_12_  (.A(\M1/stage1/carry0 [3]),
    .B(\M1/stage1/carry1 [3]),
    .S(\M1/stage1/_02_ ),
    .Z(\M1/c1 ));
 AND2_X1 \M1/stage1/gen_csa[1].FA0/HA1/_0_  (.A1(\M1/prodm1 [1]),
    .A2(\M1/prodm2 [1]),
    .ZN(\M1/stage1/gen_csa[1].FA0/ha1_carry ));
 XOR2_X2 \M1/stage1/gen_csa[1].FA0/HA1/_1_  (.A(\M1/prodm1 [1]),
    .B(\M1/prodm2 [1]),
    .Z(\M1/stage1/gen_csa[1].FA0/ha1_sum ));
 AND2_X1 \M1/stage1/gen_csa[1].FA0/HA2/_0_  (.A1(\M1/stage1/gen_csa[1].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M1/stage1/gen_csa[1].FA0/ha2_carry ));
 XOR2_X1 \M1/stage1/gen_csa[1].FA0/HA2/_1_  (.A(\M1/stage1/gen_csa[1].FA0/ha1_sum ),
    .B(ground),
    .Z(\M1/stage1/sum0 [1]));
 OR2_X1 \M1/stage1/gen_csa[1].FA0/_0_  (.A1(\M1/stage1/gen_csa[1].FA0/ha1_carry ),
    .A2(\M1/stage1/gen_csa[1].FA0/ha2_carry ),
    .ZN(\M1/stage1/carry0 [1]));
 AND2_X1 \M1/stage1/gen_csa[1].FA1/HA1/_0_  (.A1(\M1/prodm1 [1]),
    .A2(\M1/prodm2 [1]),
    .ZN(\M1/stage1/gen_csa[1].FA1/ha1_carry ));
 XOR2_X2 \M1/stage1/gen_csa[1].FA1/HA1/_1_  (.A(\M1/prodm1 [1]),
    .B(\M1/prodm2 [1]),
    .Z(\M1/stage1/gen_csa[1].FA1/ha1_sum ));
 AND2_X1 \M1/stage1/gen_csa[1].FA1/HA2/_0_  (.A1(\M1/stage1/gen_csa[1].FA1/ha1_sum ),
    .A2(\M1/stage1/_03_ ),
    .ZN(\M1/stage1/gen_csa[1].FA1/ha2_carry ));
 XOR2_X1 \M1/stage1/gen_csa[1].FA1/HA2/_1_  (.A(\M1/stage1/gen_csa[1].FA1/ha1_sum ),
    .B(\M1/stage1/_03_ ),
    .Z(\M1/stage1/sum1 [1]));
 OR2_X1 \M1/stage1/gen_csa[1].FA1/_0_  (.A1(\M1/stage1/gen_csa[1].FA1/ha1_carry ),
    .A2(\M1/stage1/gen_csa[1].FA1/ha2_carry ),
    .ZN(\M1/stage1/carry1 [1]));
 AND2_X1 \M1/stage1/gen_csa[2].FA0/HA1/_0_  (.A1(\M1/prodm1 [2]),
    .A2(\M1/prodm2 [2]),
    .ZN(\M1/stage1/gen_csa[2].FA0/ha1_carry ));
 XOR2_X1 \M1/stage1/gen_csa[2].FA0/HA1/_1_  (.A(\M1/prodm1 [2]),
    .B(\M1/prodm2 [2]),
    .Z(\M1/stage1/gen_csa[2].FA0/ha1_sum ));
 AND2_X1 \M1/stage1/gen_csa[2].FA0/HA2/_0_  (.A1(\M1/stage1/gen_csa[2].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M1/stage1/gen_csa[2].FA0/ha2_carry ));
 XOR2_X1 \M1/stage1/gen_csa[2].FA0/HA2/_1_  (.A(\M1/stage1/gen_csa[2].FA0/ha1_sum ),
    .B(ground),
    .Z(\M1/stage1/sum0 [2]));
 OR2_X1 \M1/stage1/gen_csa[2].FA0/_0_  (.A1(\M1/stage1/gen_csa[2].FA0/ha1_carry ),
    .A2(\M1/stage1/gen_csa[2].FA0/ha2_carry ),
    .ZN(\M1/stage1/carry0 [2]));
 AND2_X1 \M1/stage1/gen_csa[2].FA1/HA1/_0_  (.A1(\M1/prodm1 [2]),
    .A2(\M1/prodm2 [2]),
    .ZN(\M1/stage1/gen_csa[2].FA1/ha1_carry ));
 XOR2_X2 \M1/stage1/gen_csa[2].FA1/HA1/_1_  (.A(\M1/prodm1 [2]),
    .B(\M1/prodm2 [2]),
    .Z(\M1/stage1/gen_csa[2].FA1/ha1_sum ));
 AND2_X1 \M1/stage1/gen_csa[2].FA1/HA2/_0_  (.A1(\M1/stage1/gen_csa[2].FA1/ha1_sum ),
    .A2(\M1/stage1/_03_ ),
    .ZN(\M1/stage1/gen_csa[2].FA1/ha2_carry ));
 XOR2_X1 \M1/stage1/gen_csa[2].FA1/HA2/_1_  (.A(\M1/stage1/gen_csa[2].FA1/ha1_sum ),
    .B(\M1/stage1/_03_ ),
    .Z(\M1/stage1/sum1 [2]));
 OR2_X1 \M1/stage1/gen_csa[2].FA1/_0_  (.A1(\M1/stage1/gen_csa[2].FA1/ha1_carry ),
    .A2(\M1/stage1/gen_csa[2].FA1/ha2_carry ),
    .ZN(\M1/stage1/carry1 [2]));
 AND2_X1 \M1/stage1/gen_csa[3].FA0/HA1/_0_  (.A1(\M1/prodm1 [3]),
    .A2(\M1/prodm2 [3]),
    .ZN(\M1/stage1/gen_csa[3].FA0/ha1_carry ));
 XOR2_X2 \M1/stage1/gen_csa[3].FA0/HA1/_1_  (.A(\M1/prodm1 [3]),
    .B(\M1/prodm2 [3]),
    .Z(\M1/stage1/gen_csa[3].FA0/ha1_sum ));
 AND2_X1 \M1/stage1/gen_csa[3].FA0/HA2/_0_  (.A1(\M1/stage1/gen_csa[3].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M1/stage1/gen_csa[3].FA0/ha2_carry ));
 XOR2_X1 \M1/stage1/gen_csa[3].FA0/HA2/_1_  (.A(\M1/stage1/gen_csa[3].FA0/ha1_sum ),
    .B(ground),
    .Z(\M1/stage1/sum0 [3]));
 OR2_X1 \M1/stage1/gen_csa[3].FA0/_0_  (.A1(\M1/stage1/gen_csa[3].FA0/ha1_carry ),
    .A2(\M1/stage1/gen_csa[3].FA0/ha2_carry ),
    .ZN(\M1/stage1/carry0 [3]));
 AND2_X1 \M1/stage1/gen_csa[3].FA1/HA1/_0_  (.A1(\M1/prodm1 [3]),
    .A2(\M1/prodm2 [3]),
    .ZN(\M1/stage1/gen_csa[3].FA1/ha1_carry ));
 XOR2_X2 \M1/stage1/gen_csa[3].FA1/HA1/_1_  (.A(\M1/prodm1 [3]),
    .B(\M1/prodm2 [3]),
    .Z(\M1/stage1/gen_csa[3].FA1/ha1_sum ));
 AND2_X1 \M1/stage1/gen_csa[3].FA1/HA2/_0_  (.A1(\M1/stage1/gen_csa[3].FA1/ha1_sum ),
    .A2(\M1/stage1/_03_ ),
    .ZN(\M1/stage1/gen_csa[3].FA1/ha2_carry ));
 XOR2_X1 \M1/stage1/gen_csa[3].FA1/HA2/_1_  (.A(\M1/stage1/gen_csa[3].FA1/ha1_sum ),
    .B(\M1/stage1/_03_ ),
    .Z(\M1/stage1/sum1 [3]));
 OR2_X1 \M1/stage1/gen_csa[3].FA1/_0_  (.A1(\M1/stage1/gen_csa[3].FA1/ha1_carry ),
    .A2(\M1/stage1/gen_csa[3].FA1/ha2_carry ),
    .ZN(\M1/stage1/carry1 [3]));
 AND2_X1 \M1/stage2/FA1_0/HA1/_0_  (.A1(\M1/prodm0 [2]),
    .A2(\M1/sums1 [0]),
    .ZN(\M1/stage2/FA1_0/ha1_carry ));
 XOR2_X2 \M1/stage2/FA1_0/HA1/_1_  (.A(\M1/prodm0 [2]),
    .B(\M1/sums1 [0]),
    .Z(\M1/stage2/FA1_0/ha1_sum ));
 AND2_X1 \M1/stage2/FA1_0/HA2/_0_  (.A1(\M1/stage2/FA1_0/ha1_sum ),
    .A2(\M1/stage2/_03_ ),
    .ZN(\M1/stage2/FA1_0/ha2_carry ));
 XOR2_X1 \M1/stage2/FA1_0/HA2/_1_  (.A(\M1/stage2/FA1_0/ha1_sum ),
    .B(\M1/stage2/_03_ ),
    .Z(\M1/stage2/sum1 [0]));
 OR2_X1 \M1/stage2/FA1_0/_0_  (.A1(\M1/stage2/FA1_0/ha1_carry ),
    .A2(\M1/stage2/FA1_0/ha2_carry ),
    .ZN(\M1/stage2/carry1 [0]));
 AND2_X1 \M1/stage2/HA0_0/_0_  (.A1(\M1/prodm0 [2]),
    .A2(\M1/sums1 [0]),
    .ZN(\M1/stage2/carry0 [0]));
 XOR2_X1 \M1/stage2/HA0_0/_1_  (.A(\M1/prodm0 [2]),
    .B(\M1/sums1 [0]),
    .Z(\M1/stage2/sum0 [0]));
 INV_X2 \M1/stage2/_04_  (.A(ground),
    .ZN(\M1/stage2/_03_ ));
 MUX2_X1 \M1/stage2/_05_  (.A(\M1/stage2/sum0 [0]),
    .B(\M1/stage2/sum1 [0]),
    .S(ground),
    .Z(prodm1[2]));
 MUX2_X1 \M1/stage2/_06_  (.A(\M1/stage2/carry0 [0]),
    .B(\M1/stage2/carry1 [0]),
    .S(ground),
    .Z(\M1/stage2/_00_ ));
 MUX2_X1 \M1/stage2/_07_  (.A(\M1/stage2/sum0 [1]),
    .B(\M1/stage2/sum1 [1]),
    .S(\M1/stage2/_00_ ),
    .Z(prodm1[3]));
 MUX2_X1 \M1/stage2/_08_  (.A(\M1/stage2/carry0 [1]),
    .B(\M1/stage2/carry1 [1]),
    .S(\M1/stage2/_00_ ),
    .Z(\M1/stage2/_01_ ));
 MUX2_X2 \M1/stage2/_09_  (.A(\M1/stage2/sum0 [2]),
    .B(\M1/stage2/sum1 [2]),
    .S(\M1/stage2/_01_ ),
    .Z(\M1/sums2 [2]));
 MUX2_X1 \M1/stage2/_10_  (.A(\M1/stage2/carry0 [2]),
    .B(\M1/stage2/carry1 [2]),
    .S(\M1/stage2/_01_ ),
    .Z(\M1/stage2/_02_ ));
 MUX2_X2 \M1/stage2/_11_  (.A(\M1/stage2/sum0 [3]),
    .B(\M1/stage2/sum1 [3]),
    .S(\M1/stage2/_02_ ),
    .Z(\M1/sums2 [3]));
 MUX2_X1 \M1/stage2/_12_  (.A(\M1/stage2/carry0 [3]),
    .B(\M1/stage2/carry1 [3]),
    .S(\M1/stage2/_02_ ),
    .Z(\M1/c2 ));
 AND2_X1 \M1/stage2/gen_csa[1].FA0/HA1/_0_  (.A1(\M1/prodm0 [3]),
    .A2(\M1/sums1 [1]),
    .ZN(\M1/stage2/gen_csa[1].FA0/ha1_carry ));
 XOR2_X2 \M1/stage2/gen_csa[1].FA0/HA1/_1_  (.A(\M1/prodm0 [3]),
    .B(\M1/sums1 [1]),
    .Z(\M1/stage2/gen_csa[1].FA0/ha1_sum ));
 AND2_X1 \M1/stage2/gen_csa[1].FA0/HA2/_0_  (.A1(\M1/stage2/gen_csa[1].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M1/stage2/gen_csa[1].FA0/ha2_carry ));
 XOR2_X1 \M1/stage2/gen_csa[1].FA0/HA2/_1_  (.A(\M1/stage2/gen_csa[1].FA0/ha1_sum ),
    .B(ground),
    .Z(\M1/stage2/sum0 [1]));
 OR2_X1 \M1/stage2/gen_csa[1].FA0/_0_  (.A1(\M1/stage2/gen_csa[1].FA0/ha1_carry ),
    .A2(\M1/stage2/gen_csa[1].FA0/ha2_carry ),
    .ZN(\M1/stage2/carry0 [1]));
 AND2_X1 \M1/stage2/gen_csa[1].FA1/HA1/_0_  (.A1(\M1/prodm0 [3]),
    .A2(\M1/sums1 [1]),
    .ZN(\M1/stage2/gen_csa[1].FA1/ha1_carry ));
 XOR2_X2 \M1/stage2/gen_csa[1].FA1/HA1/_1_  (.A(\M1/prodm0 [3]),
    .B(\M1/sums1 [1]),
    .Z(\M1/stage2/gen_csa[1].FA1/ha1_sum ));
 AND2_X1 \M1/stage2/gen_csa[1].FA1/HA2/_0_  (.A1(\M1/stage2/gen_csa[1].FA1/ha1_sum ),
    .A2(\M1/stage2/_03_ ),
    .ZN(\M1/stage2/gen_csa[1].FA1/ha2_carry ));
 XOR2_X1 \M1/stage2/gen_csa[1].FA1/HA2/_1_  (.A(\M1/stage2/gen_csa[1].FA1/ha1_sum ),
    .B(\M1/stage2/_03_ ),
    .Z(\M1/stage2/sum1 [1]));
 OR2_X1 \M1/stage2/gen_csa[1].FA1/_0_  (.A1(\M1/stage2/gen_csa[1].FA1/ha1_carry ),
    .A2(\M1/stage2/gen_csa[1].FA1/ha2_carry ),
    .ZN(\M1/stage2/carry1 [1]));
 AND2_X1 \M1/stage2/gen_csa[2].FA0/HA1/_0_  (.A1(ground),
    .A2(\M1/sums1 [2]),
    .ZN(\M1/stage2/gen_csa[2].FA0/ha1_carry ));
 XOR2_X1 \M1/stage2/gen_csa[2].FA0/HA1/_1_  (.A(ground),
    .B(\M1/sums1 [2]),
    .Z(\M1/stage2/gen_csa[2].FA0/ha1_sum ));
 AND2_X1 \M1/stage2/gen_csa[2].FA0/HA2/_0_  (.A1(\M1/stage2/gen_csa[2].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M1/stage2/gen_csa[2].FA0/ha2_carry ));
 XOR2_X1 \M1/stage2/gen_csa[2].FA0/HA2/_1_  (.A(\M1/stage2/gen_csa[2].FA0/ha1_sum ),
    .B(ground),
    .Z(\M1/stage2/sum0 [2]));
 OR2_X1 \M1/stage2/gen_csa[2].FA0/_0_  (.A1(\M1/stage2/gen_csa[2].FA0/ha1_carry ),
    .A2(\M1/stage2/gen_csa[2].FA0/ha2_carry ),
    .ZN(\M1/stage2/carry0 [2]));
 AND2_X1 \M1/stage2/gen_csa[2].FA1/HA1/_0_  (.A1(ground),
    .A2(\M1/sums1 [2]),
    .ZN(\M1/stage2/gen_csa[2].FA1/ha1_carry ));
 XOR2_X2 \M1/stage2/gen_csa[2].FA1/HA1/_1_  (.A(ground),
    .B(\M1/sums1 [2]),
    .Z(\M1/stage2/gen_csa[2].FA1/ha1_sum ));
 AND2_X1 \M1/stage2/gen_csa[2].FA1/HA2/_0_  (.A1(\M1/stage2/gen_csa[2].FA1/ha1_sum ),
    .A2(\M1/stage2/_03_ ),
    .ZN(\M1/stage2/gen_csa[2].FA1/ha2_carry ));
 XOR2_X1 \M1/stage2/gen_csa[2].FA1/HA2/_1_  (.A(\M1/stage2/gen_csa[2].FA1/ha1_sum ),
    .B(\M1/stage2/_03_ ),
    .Z(\M1/stage2/sum1 [2]));
 OR2_X1 \M1/stage2/gen_csa[2].FA1/_0_  (.A1(\M1/stage2/gen_csa[2].FA1/ha1_carry ),
    .A2(\M1/stage2/gen_csa[2].FA1/ha2_carry ),
    .ZN(\M1/stage2/carry1 [2]));
 AND2_X1 \M1/stage2/gen_csa[3].FA0/HA1/_0_  (.A1(ground),
    .A2(\M1/sums1 [3]),
    .ZN(\M1/stage2/gen_csa[3].FA0/ha1_carry ));
 XOR2_X2 \M1/stage2/gen_csa[3].FA0/HA1/_1_  (.A(ground),
    .B(\M1/sums1 [3]),
    .Z(\M1/stage2/gen_csa[3].FA0/ha1_sum ));
 AND2_X1 \M1/stage2/gen_csa[3].FA0/HA2/_0_  (.A1(\M1/stage2/gen_csa[3].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M1/stage2/gen_csa[3].FA0/ha2_carry ));
 XOR2_X1 \M1/stage2/gen_csa[3].FA0/HA2/_1_  (.A(\M1/stage2/gen_csa[3].FA0/ha1_sum ),
    .B(ground),
    .Z(\M1/stage2/sum0 [3]));
 OR2_X1 \M1/stage2/gen_csa[3].FA0/_0_  (.A1(\M1/stage2/gen_csa[3].FA0/ha1_carry ),
    .A2(\M1/stage2/gen_csa[3].FA0/ha2_carry ),
    .ZN(\M1/stage2/carry0 [3]));
 AND2_X1 \M1/stage2/gen_csa[3].FA1/HA1/_0_  (.A1(ground),
    .A2(\M1/sums1 [3]),
    .ZN(\M1/stage2/gen_csa[3].FA1/ha1_carry ));
 XOR2_X2 \M1/stage2/gen_csa[3].FA1/HA1/_1_  (.A(ground),
    .B(\M1/sums1 [3]),
    .Z(\M1/stage2/gen_csa[3].FA1/ha1_sum ));
 AND2_X1 \M1/stage2/gen_csa[3].FA1/HA2/_0_  (.A1(\M1/stage2/gen_csa[3].FA1/ha1_sum ),
    .A2(\M1/stage2/_03_ ),
    .ZN(\M1/stage2/gen_csa[3].FA1/ha2_carry ));
 XOR2_X1 \M1/stage2/gen_csa[3].FA1/HA2/_1_  (.A(\M1/stage2/gen_csa[3].FA1/ha1_sum ),
    .B(\M1/stage2/_03_ ),
    .Z(\M1/stage2/sum1 [3]));
 OR2_X1 \M1/stage2/gen_csa[3].FA1/_0_  (.A1(\M1/stage2/gen_csa[3].FA1/ha1_carry ),
    .A2(\M1/stage2/gen_csa[3].FA1/ha2_carry ),
    .ZN(\M1/stage2/carry1 [3]));
 AND2_X1 \M1/stage3/FA1_0/HA1/_0_  (.A1(\M1/sums2 [2]),
    .A2(\M1/prodm3 [0]),
    .ZN(\M1/stage3/FA1_0/ha1_carry ));
 XOR2_X2 \M1/stage3/FA1_0/HA1/_1_  (.A(\M1/sums2 [2]),
    .B(\M1/prodm3 [0]),
    .Z(\M1/stage3/FA1_0/ha1_sum ));
 AND2_X1 \M1/stage3/FA1_0/HA2/_0_  (.A1(\M1/stage3/FA1_0/ha1_sum ),
    .A2(\M1/stage3/_03_ ),
    .ZN(\M1/stage3/FA1_0/ha2_carry ));
 XOR2_X1 \M1/stage3/FA1_0/HA2/_1_  (.A(\M1/stage3/FA1_0/ha1_sum ),
    .B(\M1/stage3/_03_ ),
    .Z(\M1/stage3/sum1 [0]));
 OR2_X1 \M1/stage3/FA1_0/_0_  (.A1(\M1/stage3/FA1_0/ha1_carry ),
    .A2(\M1/stage3/FA1_0/ha2_carry ),
    .ZN(\M1/stage3/carry1 [0]));
 AND2_X1 \M1/stage3/HA0_0/_0_  (.A1(\M1/sums2 [2]),
    .A2(\M1/prodm3 [0]),
    .ZN(\M1/stage3/carry0 [0]));
 XOR2_X1 \M1/stage3/HA0_0/_1_  (.A(\M1/sums2 [2]),
    .B(\M1/prodm3 [0]),
    .Z(\M1/stage3/sum0 [0]));
 INV_X2 \M1/stage3/_04_  (.A(ground),
    .ZN(\M1/stage3/_03_ ));
 MUX2_X1 \M1/stage3/_05_  (.A(\M1/stage3/sum0 [0]),
    .B(\M1/stage3/sum1 [0]),
    .S(ground),
    .Z(prodm1[4]));
 MUX2_X1 \M1/stage3/_06_  (.A(\M1/stage3/carry0 [0]),
    .B(\M1/stage3/carry1 [0]),
    .S(ground),
    .Z(\M1/stage3/_00_ ));
 MUX2_X1 \M1/stage3/_07_  (.A(\M1/stage3/sum0 [1]),
    .B(\M1/stage3/sum1 [1]),
    .S(\M1/stage3/_00_ ),
    .Z(prodm1[5]));
 MUX2_X1 \M1/stage3/_08_  (.A(\M1/stage3/carry0 [1]),
    .B(\M1/stage3/carry1 [1]),
    .S(\M1/stage3/_00_ ),
    .Z(\M1/stage3/_01_ ));
 MUX2_X1 \M1/stage3/_09_  (.A(\M1/stage3/sum0 [2]),
    .B(\M1/stage3/sum1 [2]),
    .S(\M1/stage3/_01_ ),
    .Z(prodm1[6]));
 MUX2_X1 \M1/stage3/_10_  (.A(\M1/stage3/carry0 [2]),
    .B(\M1/stage3/carry1 [2]),
    .S(\M1/stage3/_01_ ),
    .Z(\M1/stage3/_02_ ));
 MUX2_X1 \M1/stage3/_11_  (.A(\M1/stage3/sum0 [3]),
    .B(\M1/stage3/sum1 [3]),
    .S(\M1/stage3/_02_ ),
    .Z(prodm1[7]));
 MUX2_X1 \M1/stage3/_12_  (.A(\M1/stage3/carry0 [3]),
    .B(\M1/stage3/carry1 [3]),
    .S(\M1/stage3/_02_ ),
    .Z(ov2));
 AND2_X1 \M1/stage3/gen_csa[1].FA0/HA1/_0_  (.A1(\M1/sums2 [3]),
    .A2(\M1/prodm3 [1]),
    .ZN(\M1/stage3/gen_csa[1].FA0/ha1_carry ));
 XOR2_X2 \M1/stage3/gen_csa[1].FA0/HA1/_1_  (.A(\M1/sums2 [3]),
    .B(\M1/prodm3 [1]),
    .Z(\M1/stage3/gen_csa[1].FA0/ha1_sum ));
 AND2_X1 \M1/stage3/gen_csa[1].FA0/HA2/_0_  (.A1(\M1/stage3/gen_csa[1].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M1/stage3/gen_csa[1].FA0/ha2_carry ));
 XOR2_X1 \M1/stage3/gen_csa[1].FA0/HA2/_1_  (.A(\M1/stage3/gen_csa[1].FA0/ha1_sum ),
    .B(ground),
    .Z(\M1/stage3/sum0 [1]));
 OR2_X1 \M1/stage3/gen_csa[1].FA0/_0_  (.A1(\M1/stage3/gen_csa[1].FA0/ha1_carry ),
    .A2(\M1/stage3/gen_csa[1].FA0/ha2_carry ),
    .ZN(\M1/stage3/carry0 [1]));
 AND2_X1 \M1/stage3/gen_csa[1].FA1/HA1/_0_  (.A1(\M1/sums2 [3]),
    .A2(\M1/prodm3 [1]),
    .ZN(\M1/stage3/gen_csa[1].FA1/ha1_carry ));
 XOR2_X2 \M1/stage3/gen_csa[1].FA1/HA1/_1_  (.A(\M1/sums2 [3]),
    .B(\M1/prodm3 [1]),
    .Z(\M1/stage3/gen_csa[1].FA1/ha1_sum ));
 AND2_X1 \M1/stage3/gen_csa[1].FA1/HA2/_0_  (.A1(\M1/stage3/gen_csa[1].FA1/ha1_sum ),
    .A2(\M1/stage3/_03_ ),
    .ZN(\M1/stage3/gen_csa[1].FA1/ha2_carry ));
 XOR2_X1 \M1/stage3/gen_csa[1].FA1/HA2/_1_  (.A(\M1/stage3/gen_csa[1].FA1/ha1_sum ),
    .B(\M1/stage3/_03_ ),
    .Z(\M1/stage3/sum1 [1]));
 OR2_X1 \M1/stage3/gen_csa[1].FA1/_0_  (.A1(\M1/stage3/gen_csa[1].FA1/ha1_carry ),
    .A2(\M1/stage3/gen_csa[1].FA1/ha2_carry ),
    .ZN(\M1/stage3/carry1 [1]));
 AND2_X1 \M1/stage3/gen_csa[2].FA0/HA1/_0_  (.A1(\M1/cnet ),
    .A2(\M1/prodm3 [2]),
    .ZN(\M1/stage3/gen_csa[2].FA0/ha1_carry ));
 XOR2_X2 \M1/stage3/gen_csa[2].FA0/HA1/_1_  (.A(\M1/cnet ),
    .B(\M1/prodm3 [2]),
    .Z(\M1/stage3/gen_csa[2].FA0/ha1_sum ));
 AND2_X1 \M1/stage3/gen_csa[2].FA0/HA2/_0_  (.A1(\M1/stage3/gen_csa[2].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M1/stage3/gen_csa[2].FA0/ha2_carry ));
 XOR2_X1 \M1/stage3/gen_csa[2].FA0/HA2/_1_  (.A(\M1/stage3/gen_csa[2].FA0/ha1_sum ),
    .B(ground),
    .Z(\M1/stage3/sum0 [2]));
 OR2_X1 \M1/stage3/gen_csa[2].FA0/_0_  (.A1(\M1/stage3/gen_csa[2].FA0/ha1_carry ),
    .A2(\M1/stage3/gen_csa[2].FA0/ha2_carry ),
    .ZN(\M1/stage3/carry0 [2]));
 AND2_X1 \M1/stage3/gen_csa[2].FA1/HA1/_0_  (.A1(\M1/cnet ),
    .A2(\M1/prodm3 [2]),
    .ZN(\M1/stage3/gen_csa[2].FA1/ha1_carry ));
 XOR2_X2 \M1/stage3/gen_csa[2].FA1/HA1/_1_  (.A(\M1/cnet ),
    .B(\M1/prodm3 [2]),
    .Z(\M1/stage3/gen_csa[2].FA1/ha1_sum ));
 AND2_X1 \M1/stage3/gen_csa[2].FA1/HA2/_0_  (.A1(\M1/stage3/gen_csa[2].FA1/ha1_sum ),
    .A2(\M1/stage3/_03_ ),
    .ZN(\M1/stage3/gen_csa[2].FA1/ha2_carry ));
 XOR2_X1 \M1/stage3/gen_csa[2].FA1/HA2/_1_  (.A(\M1/stage3/gen_csa[2].FA1/ha1_sum ),
    .B(\M1/stage3/_03_ ),
    .Z(\M1/stage3/sum1 [2]));
 OR2_X1 \M1/stage3/gen_csa[2].FA1/_0_  (.A1(\M1/stage3/gen_csa[2].FA1/ha1_carry ),
    .A2(\M1/stage3/gen_csa[2].FA1/ha2_carry ),
    .ZN(\M1/stage3/carry1 [2]));
 AND2_X1 \M1/stage3/gen_csa[3].FA0/HA1/_0_  (.A1(ground),
    .A2(\M1/prodm3 [3]),
    .ZN(\M1/stage3/gen_csa[3].FA0/ha1_carry ));
 XOR2_X1 \M1/stage3/gen_csa[3].FA0/HA1/_1_  (.A(ground),
    .B(\M1/prodm3 [3]),
    .Z(\M1/stage3/gen_csa[3].FA0/ha1_sum ));
 AND2_X1 \M1/stage3/gen_csa[3].FA0/HA2/_0_  (.A1(\M1/stage3/gen_csa[3].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M1/stage3/gen_csa[3].FA0/ha2_carry ));
 XOR2_X1 \M1/stage3/gen_csa[3].FA0/HA2/_1_  (.A(\M1/stage3/gen_csa[3].FA0/ha1_sum ),
    .B(ground),
    .Z(\M1/stage3/sum0 [3]));
 OR2_X1 \M1/stage3/gen_csa[3].FA0/_0_  (.A1(\M1/stage3/gen_csa[3].FA0/ha1_carry ),
    .A2(\M1/stage3/gen_csa[3].FA0/ha2_carry ),
    .ZN(\M1/stage3/carry0 [3]));
 AND2_X1 \M1/stage3/gen_csa[3].FA1/HA1/_0_  (.A1(ground),
    .A2(\M1/prodm3 [3]),
    .ZN(\M1/stage3/gen_csa[3].FA1/ha1_carry ));
 XOR2_X2 \M1/stage3/gen_csa[3].FA1/HA1/_1_  (.A(ground),
    .B(\M1/prodm3 [3]),
    .Z(\M1/stage3/gen_csa[3].FA1/ha1_sum ));
 AND2_X1 \M1/stage3/gen_csa[3].FA1/HA2/_0_  (.A1(\M1/stage3/gen_csa[3].FA1/ha1_sum ),
    .A2(\M1/stage3/_03_ ),
    .ZN(\M1/stage3/gen_csa[3].FA1/ha2_carry ));
 XOR2_X1 \M1/stage3/gen_csa[3].FA1/HA2/_1_  (.A(\M1/stage3/gen_csa[3].FA1/ha1_sum ),
    .B(\M1/stage3/_03_ ),
    .Z(\M1/stage3/sum1 [3]));
 OR2_X1 \M1/stage3/gen_csa[3].FA1/_0_  (.A1(\M1/stage3/gen_csa[3].FA1/ha1_carry ),
    .A2(\M1/stage3/gen_csa[3].FA1/ha2_carry ),
    .ZN(\M1/stage3/carry1 [3]));
 AND2_X1 \M2/M0/HA0/_0_  (.A1(\M2/M0/a0b1 ),
    .A2(\M2/M0/a1b0 ),
    .ZN(\M2/M0/carry ));
 XOR2_X1 \M2/M0/HA0/_1_  (.A(\M2/M0/a0b1 ),
    .B(\M2/M0/a1b0 ),
    .Z(prodm2[1]));
 AND2_X1 \M2/M0/HA1/_0_  (.A1(\M2/M0/a1b1 ),
    .A2(\M2/M0/carry ),
    .ZN(\M2/prodm0 [3]));
 XOR2_X2 \M2/M0/HA1/_1_  (.A(\M2/M0/a1b1 ),
    .B(\M2/M0/carry ),
    .Z(\M2/prodm0 [2]));
 AND2_X1 \M2/M0/_0_  (.A1(a[5]),
    .A2(b[1]),
    .ZN(\M2/M0/a1b1 ));
 AND2_X1 \M2/M0/_1_  (.A1(b[1]),
    .A2(a[4]),
    .ZN(\M2/M0/a0b1 ));
 AND2_X1 \M2/M0/_2_  (.A1(a[5]),
    .A2(b[0]),
    .ZN(\M2/M0/a1b0 ));
 AND2_X1 \M2/M0/_3_  (.A1(a[4]),
    .A2(b[0]),
    .ZN(prodm2[0]));
 AND2_X1 \M2/M1/HA0/_0_  (.A1(\M2/M1/a0b1 ),
    .A2(\M2/M1/a1b0 ),
    .ZN(\M2/M1/carry ));
 XOR2_X2 \M2/M1/HA0/_1_  (.A(\M2/M1/a0b1 ),
    .B(\M2/M1/a1b0 ),
    .Z(\M2/prodm1 [1]));
 AND2_X1 \M2/M1/HA1/_0_  (.A1(\M2/M1/a1b1 ),
    .A2(\M2/M1/carry ),
    .ZN(\M2/prodm1 [3]));
 XOR2_X2 \M2/M1/HA1/_1_  (.A(\M2/M1/a1b1 ),
    .B(\M2/M1/carry ),
    .Z(\M2/prodm1 [2]));
 AND2_X1 \M2/M1/_0_  (.A1(a[5]),
    .A2(b[3]),
    .ZN(\M2/M1/a1b1 ));
 AND2_X1 \M2/M1/_1_  (.A1(b[3]),
    .A2(a[4]),
    .ZN(\M2/M1/a0b1 ));
 AND2_X1 \M2/M1/_2_  (.A1(a[5]),
    .A2(b[2]),
    .ZN(\M2/M1/a1b0 ));
 AND2_X1 \M2/M1/_3_  (.A1(a[4]),
    .A2(b[2]),
    .ZN(\M2/prodm1 [0]));
 AND2_X1 \M2/M2/HA0/_0_  (.A1(\M2/M2/a0b1 ),
    .A2(\M2/M2/a1b0 ),
    .ZN(\M2/M2/carry ));
 XOR2_X2 \M2/M2/HA0/_1_  (.A(\M2/M2/a0b1 ),
    .B(\M2/M2/a1b0 ),
    .Z(\M2/prodm2 [1]));
 AND2_X1 \M2/M2/HA1/_0_  (.A1(\M2/M2/a1b1 ),
    .A2(\M2/M2/carry ),
    .ZN(\M2/prodm2 [3]));
 XOR2_X2 \M2/M2/HA1/_1_  (.A(\M2/M2/a1b1 ),
    .B(\M2/M2/carry ),
    .Z(\M2/prodm2 [2]));
 AND2_X1 \M2/M2/_0_  (.A1(a[7]),
    .A2(b[1]),
    .ZN(\M2/M2/a1b1 ));
 AND2_X1 \M2/M2/_1_  (.A1(b[1]),
    .A2(a[6]),
    .ZN(\M2/M2/a0b1 ));
 AND2_X1 \M2/M2/_2_  (.A1(a[7]),
    .A2(b[0]),
    .ZN(\M2/M2/a1b0 ));
 AND2_X1 \M2/M2/_3_  (.A1(a[6]),
    .A2(b[0]),
    .ZN(\M2/prodm2 [0]));
 AND2_X1 \M2/M3/HA0/_0_  (.A1(\M2/M3/a0b1 ),
    .A2(\M2/M3/a1b0 ),
    .ZN(\M2/M3/carry ));
 XOR2_X2 \M2/M3/HA0/_1_  (.A(\M2/M3/a0b1 ),
    .B(\M2/M3/a1b0 ),
    .Z(\M2/prodm3 [1]));
 AND2_X2 \M2/M3/HA1/_0_  (.A1(\M2/M3/a1b1 ),
    .A2(\M2/M3/carry ),
    .ZN(\M2/prodm3 [3]));
 XOR2_X2 \M2/M3/HA1/_1_  (.A(\M2/M3/a1b1 ),
    .B(\M2/M3/carry ),
    .Z(\M2/prodm3 [2]));
 AND2_X1 \M2/M3/_0_  (.A1(a[7]),
    .A2(b[3]),
    .ZN(\M2/M3/a1b1 ));
 AND2_X1 \M2/M3/_1_  (.A1(b[3]),
    .A2(a[6]),
    .ZN(\M2/M3/a0b1 ));
 AND2_X1 \M2/M3/_2_  (.A1(a[7]),
    .A2(b[2]),
    .ZN(\M2/M3/a1b0 ));
 AND2_X1 \M2/M3/_3_  (.A1(a[6]),
    .A2(b[2]),
    .ZN(\M2/prodm3 [0]));
 OR2_X2 \M2/_0_  (.A1(\M2/c1 ),
    .A2(\M2/c2 ),
    .ZN(\M2/cnet ));
 AND2_X1 \M2/stage1/FA1_0/HA1/_0_  (.A1(\M2/prodm1 [0]),
    .A2(\M2/prodm2 [0]),
    .ZN(\M2/stage1/FA1_0/ha1_carry ));
 XOR2_X1 \M2/stage1/FA1_0/HA1/_1_  (.A(\M2/prodm1 [0]),
    .B(\M2/prodm2 [0]),
    .Z(\M2/stage1/FA1_0/ha1_sum ));
 AND2_X1 \M2/stage1/FA1_0/HA2/_0_  (.A1(\M2/stage1/FA1_0/ha1_sum ),
    .A2(\M2/stage1/_03_ ),
    .ZN(\M2/stage1/FA1_0/ha2_carry ));
 XOR2_X1 \M2/stage1/FA1_0/HA2/_1_  (.A(\M2/stage1/FA1_0/ha1_sum ),
    .B(\M2/stage1/_03_ ),
    .Z(\M2/stage1/sum1 [0]));
 OR2_X1 \M2/stage1/FA1_0/_0_  (.A1(\M2/stage1/FA1_0/ha1_carry ),
    .A2(\M2/stage1/FA1_0/ha2_carry ),
    .ZN(\M2/stage1/carry1 [0]));
 AND2_X1 \M2/stage1/HA0_0/_0_  (.A1(\M2/prodm1 [0]),
    .A2(\M2/prodm2 [0]),
    .ZN(\M2/stage1/carry0 [0]));
 XOR2_X1 \M2/stage1/HA0_0/_1_  (.A(\M2/prodm1 [0]),
    .B(\M2/prodm2 [0]),
    .Z(\M2/stage1/sum0 [0]));
 INV_X2 \M2/stage1/_04_  (.A(ground),
    .ZN(\M2/stage1/_03_ ));
 MUX2_X2 \M2/stage1/_05_  (.A(\M2/stage1/sum0 [0]),
    .B(\M2/stage1/sum1 [0]),
    .S(ground),
    .Z(\M2/sums1 [0]));
 MUX2_X1 \M2/stage1/_06_  (.A(\M2/stage1/carry0 [0]),
    .B(\M2/stage1/carry1 [0]),
    .S(ground),
    .Z(\M2/stage1/_00_ ));
 MUX2_X2 \M2/stage1/_07_  (.A(\M2/stage1/sum0 [1]),
    .B(\M2/stage1/sum1 [1]),
    .S(\M2/stage1/_00_ ),
    .Z(\M2/sums1 [1]));
 MUX2_X1 \M2/stage1/_08_  (.A(\M2/stage1/carry0 [1]),
    .B(\M2/stage1/carry1 [1]),
    .S(\M2/stage1/_00_ ),
    .Z(\M2/stage1/_01_ ));
 MUX2_X2 \M2/stage1/_09_  (.A(\M2/stage1/sum0 [2]),
    .B(\M2/stage1/sum1 [2]),
    .S(\M2/stage1/_01_ ),
    .Z(\M2/sums1 [2]));
 MUX2_X1 \M2/stage1/_10_  (.A(\M2/stage1/carry0 [2]),
    .B(\M2/stage1/carry1 [2]),
    .S(\M2/stage1/_01_ ),
    .Z(\M2/stage1/_02_ ));
 MUX2_X2 \M2/stage1/_11_  (.A(\M2/stage1/sum0 [3]),
    .B(\M2/stage1/sum1 [3]),
    .S(\M2/stage1/_02_ ),
    .Z(\M2/sums1 [3]));
 MUX2_X1 \M2/stage1/_12_  (.A(\M2/stage1/carry0 [3]),
    .B(\M2/stage1/carry1 [3]),
    .S(\M2/stage1/_02_ ),
    .Z(\M2/c1 ));
 AND2_X1 \M2/stage1/gen_csa[1].FA0/HA1/_0_  (.A1(\M2/prodm1 [1]),
    .A2(\M2/prodm2 [1]),
    .ZN(\M2/stage1/gen_csa[1].FA0/ha1_carry ));
 XOR2_X2 \M2/stage1/gen_csa[1].FA0/HA1/_1_  (.A(\M2/prodm1 [1]),
    .B(\M2/prodm2 [1]),
    .Z(\M2/stage1/gen_csa[1].FA0/ha1_sum ));
 AND2_X1 \M2/stage1/gen_csa[1].FA0/HA2/_0_  (.A1(\M2/stage1/gen_csa[1].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M2/stage1/gen_csa[1].FA0/ha2_carry ));
 XOR2_X1 \M2/stage1/gen_csa[1].FA0/HA2/_1_  (.A(\M2/stage1/gen_csa[1].FA0/ha1_sum ),
    .B(ground),
    .Z(\M2/stage1/sum0 [1]));
 OR2_X1 \M2/stage1/gen_csa[1].FA0/_0_  (.A1(\M2/stage1/gen_csa[1].FA0/ha1_carry ),
    .A2(\M2/stage1/gen_csa[1].FA0/ha2_carry ),
    .ZN(\M2/stage1/carry0 [1]));
 AND2_X1 \M2/stage1/gen_csa[1].FA1/HA1/_0_  (.A1(\M2/prodm1 [1]),
    .A2(\M2/prodm2 [1]),
    .ZN(\M2/stage1/gen_csa[1].FA1/ha1_carry ));
 XOR2_X2 \M2/stage1/gen_csa[1].FA1/HA1/_1_  (.A(\M2/prodm1 [1]),
    .B(\M2/prodm2 [1]),
    .Z(\M2/stage1/gen_csa[1].FA1/ha1_sum ));
 AND2_X1 \M2/stage1/gen_csa[1].FA1/HA2/_0_  (.A1(\M2/stage1/gen_csa[1].FA1/ha1_sum ),
    .A2(\M2/stage1/_03_ ),
    .ZN(\M2/stage1/gen_csa[1].FA1/ha2_carry ));
 XOR2_X1 \M2/stage1/gen_csa[1].FA1/HA2/_1_  (.A(\M2/stage1/gen_csa[1].FA1/ha1_sum ),
    .B(\M2/stage1/_03_ ),
    .Z(\M2/stage1/sum1 [1]));
 OR2_X1 \M2/stage1/gen_csa[1].FA1/_0_  (.A1(\M2/stage1/gen_csa[1].FA1/ha1_carry ),
    .A2(\M2/stage1/gen_csa[1].FA1/ha2_carry ),
    .ZN(\M2/stage1/carry1 [1]));
 AND2_X1 \M2/stage1/gen_csa[2].FA0/HA1/_0_  (.A1(\M2/prodm1 [2]),
    .A2(\M2/prodm2 [2]),
    .ZN(\M2/stage1/gen_csa[2].FA0/ha1_carry ));
 XOR2_X2 \M2/stage1/gen_csa[2].FA0/HA1/_1_  (.A(\M2/prodm1 [2]),
    .B(\M2/prodm2 [2]),
    .Z(\M2/stage1/gen_csa[2].FA0/ha1_sum ));
 AND2_X1 \M2/stage1/gen_csa[2].FA0/HA2/_0_  (.A1(\M2/stage1/gen_csa[2].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M2/stage1/gen_csa[2].FA0/ha2_carry ));
 XOR2_X1 \M2/stage1/gen_csa[2].FA0/HA2/_1_  (.A(\M2/stage1/gen_csa[2].FA0/ha1_sum ),
    .B(ground),
    .Z(\M2/stage1/sum0 [2]));
 OR2_X1 \M2/stage1/gen_csa[2].FA0/_0_  (.A1(\M2/stage1/gen_csa[2].FA0/ha1_carry ),
    .A2(\M2/stage1/gen_csa[2].FA0/ha2_carry ),
    .ZN(\M2/stage1/carry0 [2]));
 AND2_X1 \M2/stage1/gen_csa[2].FA1/HA1/_0_  (.A1(\M2/prodm1 [2]),
    .A2(\M2/prodm2 [2]),
    .ZN(\M2/stage1/gen_csa[2].FA1/ha1_carry ));
 XOR2_X2 \M2/stage1/gen_csa[2].FA1/HA1/_1_  (.A(\M2/prodm1 [2]),
    .B(\M2/prodm2 [2]),
    .Z(\M2/stage1/gen_csa[2].FA1/ha1_sum ));
 AND2_X1 \M2/stage1/gen_csa[2].FA1/HA2/_0_  (.A1(\M2/stage1/gen_csa[2].FA1/ha1_sum ),
    .A2(\M2/stage1/_03_ ),
    .ZN(\M2/stage1/gen_csa[2].FA1/ha2_carry ));
 XOR2_X1 \M2/stage1/gen_csa[2].FA1/HA2/_1_  (.A(\M2/stage1/gen_csa[2].FA1/ha1_sum ),
    .B(\M2/stage1/_03_ ),
    .Z(\M2/stage1/sum1 [2]));
 OR2_X1 \M2/stage1/gen_csa[2].FA1/_0_  (.A1(\M2/stage1/gen_csa[2].FA1/ha1_carry ),
    .A2(\M2/stage1/gen_csa[2].FA1/ha2_carry ),
    .ZN(\M2/stage1/carry1 [2]));
 AND2_X1 \M2/stage1/gen_csa[3].FA0/HA1/_0_  (.A1(\M2/prodm1 [3]),
    .A2(\M2/prodm2 [3]),
    .ZN(\M2/stage1/gen_csa[3].FA0/ha1_carry ));
 XOR2_X1 \M2/stage1/gen_csa[3].FA0/HA1/_1_  (.A(\M2/prodm1 [3]),
    .B(\M2/prodm2 [3]),
    .Z(\M2/stage1/gen_csa[3].FA0/ha1_sum ));
 AND2_X1 \M2/stage1/gen_csa[3].FA0/HA2/_0_  (.A1(\M2/stage1/gen_csa[3].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M2/stage1/gen_csa[3].FA0/ha2_carry ));
 XOR2_X1 \M2/stage1/gen_csa[3].FA0/HA2/_1_  (.A(\M2/stage1/gen_csa[3].FA0/ha1_sum ),
    .B(ground),
    .Z(\M2/stage1/sum0 [3]));
 OR2_X1 \M2/stage1/gen_csa[3].FA0/_0_  (.A1(\M2/stage1/gen_csa[3].FA0/ha1_carry ),
    .A2(\M2/stage1/gen_csa[3].FA0/ha2_carry ),
    .ZN(\M2/stage1/carry0 [3]));
 AND2_X1 \M2/stage1/gen_csa[3].FA1/HA1/_0_  (.A1(\M2/prodm1 [3]),
    .A2(\M2/prodm2 [3]),
    .ZN(\M2/stage1/gen_csa[3].FA1/ha1_carry ));
 XOR2_X2 \M2/stage1/gen_csa[3].FA1/HA1/_1_  (.A(\M2/prodm1 [3]),
    .B(\M2/prodm2 [3]),
    .Z(\M2/stage1/gen_csa[3].FA1/ha1_sum ));
 AND2_X1 \M2/stage1/gen_csa[3].FA1/HA2/_0_  (.A1(\M2/stage1/gen_csa[3].FA1/ha1_sum ),
    .A2(\M2/stage1/_03_ ),
    .ZN(\M2/stage1/gen_csa[3].FA1/ha2_carry ));
 XOR2_X1 \M2/stage1/gen_csa[3].FA1/HA2/_1_  (.A(\M2/stage1/gen_csa[3].FA1/ha1_sum ),
    .B(\M2/stage1/_03_ ),
    .Z(\M2/stage1/sum1 [3]));
 OR2_X1 \M2/stage1/gen_csa[3].FA1/_0_  (.A1(\M2/stage1/gen_csa[3].FA1/ha1_carry ),
    .A2(\M2/stage1/gen_csa[3].FA1/ha2_carry ),
    .ZN(\M2/stage1/carry1 [3]));
 AND2_X1 \M2/stage2/FA1_0/HA1/_0_  (.A1(\M2/prodm0 [2]),
    .A2(\M2/sums1 [0]),
    .ZN(\M2/stage2/FA1_0/ha1_carry ));
 XOR2_X2 \M2/stage2/FA1_0/HA1/_1_  (.A(\M2/prodm0 [2]),
    .B(\M2/sums1 [0]),
    .Z(\M2/stage2/FA1_0/ha1_sum ));
 AND2_X1 \M2/stage2/FA1_0/HA2/_0_  (.A1(\M2/stage2/FA1_0/ha1_sum ),
    .A2(\M2/stage2/_03_ ),
    .ZN(\M2/stage2/FA1_0/ha2_carry ));
 XOR2_X1 \M2/stage2/FA1_0/HA2/_1_  (.A(\M2/stage2/FA1_0/ha1_sum ),
    .B(\M2/stage2/_03_ ),
    .Z(\M2/stage2/sum1 [0]));
 OR2_X1 \M2/stage2/FA1_0/_0_  (.A1(\M2/stage2/FA1_0/ha1_carry ),
    .A2(\M2/stage2/FA1_0/ha2_carry ),
    .ZN(\M2/stage2/carry1 [0]));
 AND2_X1 \M2/stage2/HA0_0/_0_  (.A1(\M2/prodm0 [2]),
    .A2(\M2/sums1 [0]),
    .ZN(\M2/stage2/carry0 [0]));
 XOR2_X1 \M2/stage2/HA0_0/_1_  (.A(\M2/prodm0 [2]),
    .B(\M2/sums1 [0]),
    .Z(\M2/stage2/sum0 [0]));
 INV_X2 \M2/stage2/_04_  (.A(ground),
    .ZN(\M2/stage2/_03_ ));
 MUX2_X1 \M2/stage2/_05_  (.A(\M2/stage2/sum0 [0]),
    .B(\M2/stage2/sum1 [0]),
    .S(ground),
    .Z(prodm2[2]));
 MUX2_X1 \M2/stage2/_06_  (.A(\M2/stage2/carry0 [0]),
    .B(\M2/stage2/carry1 [0]),
    .S(ground),
    .Z(\M2/stage2/_00_ ));
 MUX2_X1 \M2/stage2/_07_  (.A(\M2/stage2/sum0 [1]),
    .B(\M2/stage2/sum1 [1]),
    .S(\M2/stage2/_00_ ),
    .Z(prodm2[3]));
 MUX2_X1 \M2/stage2/_08_  (.A(\M2/stage2/carry0 [1]),
    .B(\M2/stage2/carry1 [1]),
    .S(\M2/stage2/_00_ ),
    .Z(\M2/stage2/_01_ ));
 MUX2_X2 \M2/stage2/_09_  (.A(\M2/stage2/sum0 [2]),
    .B(\M2/stage2/sum1 [2]),
    .S(\M2/stage2/_01_ ),
    .Z(\M2/sums2 [2]));
 MUX2_X1 \M2/stage2/_10_  (.A(\M2/stage2/carry0 [2]),
    .B(\M2/stage2/carry1 [2]),
    .S(\M2/stage2/_01_ ),
    .Z(\M2/stage2/_02_ ));
 MUX2_X2 \M2/stage2/_11_  (.A(\M2/stage2/sum0 [3]),
    .B(\M2/stage2/sum1 [3]),
    .S(\M2/stage2/_02_ ),
    .Z(\M2/sums2 [3]));
 MUX2_X1 \M2/stage2/_12_  (.A(\M2/stage2/carry0 [3]),
    .B(\M2/stage2/carry1 [3]),
    .S(\M2/stage2/_02_ ),
    .Z(\M2/c2 ));
 AND2_X1 \M2/stage2/gen_csa[1].FA0/HA1/_0_  (.A1(\M2/prodm0 [3]),
    .A2(\M2/sums1 [1]),
    .ZN(\M2/stage2/gen_csa[1].FA0/ha1_carry ));
 XOR2_X2 \M2/stage2/gen_csa[1].FA0/HA1/_1_  (.A(\M2/prodm0 [3]),
    .B(\M2/sums1 [1]),
    .Z(\M2/stage2/gen_csa[1].FA0/ha1_sum ));
 AND2_X1 \M2/stage2/gen_csa[1].FA0/HA2/_0_  (.A1(\M2/stage2/gen_csa[1].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M2/stage2/gen_csa[1].FA0/ha2_carry ));
 XOR2_X1 \M2/stage2/gen_csa[1].FA0/HA2/_1_  (.A(\M2/stage2/gen_csa[1].FA0/ha1_sum ),
    .B(ground),
    .Z(\M2/stage2/sum0 [1]));
 OR2_X1 \M2/stage2/gen_csa[1].FA0/_0_  (.A1(\M2/stage2/gen_csa[1].FA0/ha1_carry ),
    .A2(\M2/stage2/gen_csa[1].FA0/ha2_carry ),
    .ZN(\M2/stage2/carry0 [1]));
 AND2_X1 \M2/stage2/gen_csa[1].FA1/HA1/_0_  (.A1(\M2/prodm0 [3]),
    .A2(\M2/sums1 [1]),
    .ZN(\M2/stage2/gen_csa[1].FA1/ha1_carry ));
 XOR2_X2 \M2/stage2/gen_csa[1].FA1/HA1/_1_  (.A(\M2/prodm0 [3]),
    .B(\M2/sums1 [1]),
    .Z(\M2/stage2/gen_csa[1].FA1/ha1_sum ));
 AND2_X1 \M2/stage2/gen_csa[1].FA1/HA2/_0_  (.A1(\M2/stage2/gen_csa[1].FA1/ha1_sum ),
    .A2(\M2/stage2/_03_ ),
    .ZN(\M2/stage2/gen_csa[1].FA1/ha2_carry ));
 XOR2_X1 \M2/stage2/gen_csa[1].FA1/HA2/_1_  (.A(\M2/stage2/gen_csa[1].FA1/ha1_sum ),
    .B(\M2/stage2/_03_ ),
    .Z(\M2/stage2/sum1 [1]));
 OR2_X1 \M2/stage2/gen_csa[1].FA1/_0_  (.A1(\M2/stage2/gen_csa[1].FA1/ha1_carry ),
    .A2(\M2/stage2/gen_csa[1].FA1/ha2_carry ),
    .ZN(\M2/stage2/carry1 [1]));
 AND2_X1 \M2/stage2/gen_csa[2].FA0/HA1/_0_  (.A1(ground),
    .A2(\M2/sums1 [2]),
    .ZN(\M2/stage2/gen_csa[2].FA0/ha1_carry ));
 XOR2_X2 \M2/stage2/gen_csa[2].FA0/HA1/_1_  (.A(ground),
    .B(\M2/sums1 [2]),
    .Z(\M2/stage2/gen_csa[2].FA0/ha1_sum ));
 AND2_X1 \M2/stage2/gen_csa[2].FA0/HA2/_0_  (.A1(\M2/stage2/gen_csa[2].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M2/stage2/gen_csa[2].FA0/ha2_carry ));
 XOR2_X1 \M2/stage2/gen_csa[2].FA0/HA2/_1_  (.A(\M2/stage2/gen_csa[2].FA0/ha1_sum ),
    .B(ground),
    .Z(\M2/stage2/sum0 [2]));
 OR2_X1 \M2/stage2/gen_csa[2].FA0/_0_  (.A1(\M2/stage2/gen_csa[2].FA0/ha1_carry ),
    .A2(\M2/stage2/gen_csa[2].FA0/ha2_carry ),
    .ZN(\M2/stage2/carry0 [2]));
 AND2_X1 \M2/stage2/gen_csa[2].FA1/HA1/_0_  (.A1(ground),
    .A2(\M2/sums1 [2]),
    .ZN(\M2/stage2/gen_csa[2].FA1/ha1_carry ));
 XOR2_X2 \M2/stage2/gen_csa[2].FA1/HA1/_1_  (.A(ground),
    .B(\M2/sums1 [2]),
    .Z(\M2/stage2/gen_csa[2].FA1/ha1_sum ));
 AND2_X1 \M2/stage2/gen_csa[2].FA1/HA2/_0_  (.A1(\M2/stage2/gen_csa[2].FA1/ha1_sum ),
    .A2(\M2/stage2/_03_ ),
    .ZN(\M2/stage2/gen_csa[2].FA1/ha2_carry ));
 XOR2_X1 \M2/stage2/gen_csa[2].FA1/HA2/_1_  (.A(\M2/stage2/gen_csa[2].FA1/ha1_sum ),
    .B(\M2/stage2/_03_ ),
    .Z(\M2/stage2/sum1 [2]));
 OR2_X1 \M2/stage2/gen_csa[2].FA1/_0_  (.A1(\M2/stage2/gen_csa[2].FA1/ha1_carry ),
    .A2(\M2/stage2/gen_csa[2].FA1/ha2_carry ),
    .ZN(\M2/stage2/carry1 [2]));
 AND2_X1 \M2/stage2/gen_csa[3].FA0/HA1/_0_  (.A1(ground),
    .A2(\M2/sums1 [3]),
    .ZN(\M2/stage2/gen_csa[3].FA0/ha1_carry ));
 XOR2_X2 \M2/stage2/gen_csa[3].FA0/HA1/_1_  (.A(ground),
    .B(\M2/sums1 [3]),
    .Z(\M2/stage2/gen_csa[3].FA0/ha1_sum ));
 AND2_X1 \M2/stage2/gen_csa[3].FA0/HA2/_0_  (.A1(\M2/stage2/gen_csa[3].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M2/stage2/gen_csa[3].FA0/ha2_carry ));
 XOR2_X1 \M2/stage2/gen_csa[3].FA0/HA2/_1_  (.A(\M2/stage2/gen_csa[3].FA0/ha1_sum ),
    .B(ground),
    .Z(\M2/stage2/sum0 [3]));
 OR2_X1 \M2/stage2/gen_csa[3].FA0/_0_  (.A1(\M2/stage2/gen_csa[3].FA0/ha1_carry ),
    .A2(\M2/stage2/gen_csa[3].FA0/ha2_carry ),
    .ZN(\M2/stage2/carry0 [3]));
 AND2_X1 \M2/stage2/gen_csa[3].FA1/HA1/_0_  (.A1(ground),
    .A2(\M2/sums1 [3]),
    .ZN(\M2/stage2/gen_csa[3].FA1/ha1_carry ));
 XOR2_X2 \M2/stage2/gen_csa[3].FA1/HA1/_1_  (.A(ground),
    .B(\M2/sums1 [3]),
    .Z(\M2/stage2/gen_csa[3].FA1/ha1_sum ));
 AND2_X1 \M2/stage2/gen_csa[3].FA1/HA2/_0_  (.A1(\M2/stage2/gen_csa[3].FA1/ha1_sum ),
    .A2(\M2/stage2/_03_ ),
    .ZN(\M2/stage2/gen_csa[3].FA1/ha2_carry ));
 XOR2_X1 \M2/stage2/gen_csa[3].FA1/HA2/_1_  (.A(\M2/stage2/gen_csa[3].FA1/ha1_sum ),
    .B(\M2/stage2/_03_ ),
    .Z(\M2/stage2/sum1 [3]));
 OR2_X1 \M2/stage2/gen_csa[3].FA1/_0_  (.A1(\M2/stage2/gen_csa[3].FA1/ha1_carry ),
    .A2(\M2/stage2/gen_csa[3].FA1/ha2_carry ),
    .ZN(\M2/stage2/carry1 [3]));
 AND2_X1 \M2/stage3/FA1_0/HA1/_0_  (.A1(\M2/sums2 [2]),
    .A2(\M2/prodm3 [0]),
    .ZN(\M2/stage3/FA1_0/ha1_carry ));
 XOR2_X2 \M2/stage3/FA1_0/HA1/_1_  (.A(\M2/sums2 [2]),
    .B(\M2/prodm3 [0]),
    .Z(\M2/stage3/FA1_0/ha1_sum ));
 AND2_X1 \M2/stage3/FA1_0/HA2/_0_  (.A1(\M2/stage3/FA1_0/ha1_sum ),
    .A2(\M2/stage3/_03_ ),
    .ZN(\M2/stage3/FA1_0/ha2_carry ));
 XOR2_X1 \M2/stage3/FA1_0/HA2/_1_  (.A(\M2/stage3/FA1_0/ha1_sum ),
    .B(\M2/stage3/_03_ ),
    .Z(\M2/stage3/sum1 [0]));
 OR2_X1 \M2/stage3/FA1_0/_0_  (.A1(\M2/stage3/FA1_0/ha1_carry ),
    .A2(\M2/stage3/FA1_0/ha2_carry ),
    .ZN(\M2/stage3/carry1 [0]));
 AND2_X1 \M2/stage3/HA0_0/_0_  (.A1(\M2/sums2 [2]),
    .A2(\M2/prodm3 [0]),
    .ZN(\M2/stage3/carry0 [0]));
 XOR2_X1 \M2/stage3/HA0_0/_1_  (.A(\M2/sums2 [2]),
    .B(\M2/prodm3 [0]),
    .Z(\M2/stage3/sum0 [0]));
 INV_X2 \M2/stage3/_04_  (.A(ground),
    .ZN(\M2/stage3/_03_ ));
 MUX2_X1 \M2/stage3/_05_  (.A(\M2/stage3/sum0 [0]),
    .B(\M2/stage3/sum1 [0]),
    .S(ground),
    .Z(prodm2[4]));
 MUX2_X1 \M2/stage3/_06_  (.A(\M2/stage3/carry0 [0]),
    .B(\M2/stage3/carry1 [0]),
    .S(ground),
    .Z(\M2/stage3/_00_ ));
 MUX2_X1 \M2/stage3/_07_  (.A(\M2/stage3/sum0 [1]),
    .B(\M2/stage3/sum1 [1]),
    .S(\M2/stage3/_00_ ),
    .Z(prodm2[5]));
 MUX2_X1 \M2/stage3/_08_  (.A(\M2/stage3/carry0 [1]),
    .B(\M2/stage3/carry1 [1]),
    .S(\M2/stage3/_00_ ),
    .Z(\M2/stage3/_01_ ));
 MUX2_X1 \M2/stage3/_09_  (.A(\M2/stage3/sum0 [2]),
    .B(\M2/stage3/sum1 [2]),
    .S(\M2/stage3/_01_ ),
    .Z(prodm2[6]));
 MUX2_X1 \M2/stage3/_10_  (.A(\M2/stage3/carry0 [2]),
    .B(\M2/stage3/carry1 [2]),
    .S(\M2/stage3/_01_ ),
    .Z(\M2/stage3/_02_ ));
 MUX2_X1 \M2/stage3/_11_  (.A(\M2/stage3/sum0 [3]),
    .B(\M2/stage3/sum1 [3]),
    .S(\M2/stage3/_02_ ),
    .Z(prodm2[7]));
 MUX2_X1 \M2/stage3/_12_  (.A(\M2/stage3/carry0 [3]),
    .B(\M2/stage3/carry1 [3]),
    .S(\M2/stage3/_02_ ),
    .Z(ov3));
 AND2_X1 \M2/stage3/gen_csa[1].FA0/HA1/_0_  (.A1(\M2/sums2 [3]),
    .A2(\M2/prodm3 [1]),
    .ZN(\M2/stage3/gen_csa[1].FA0/ha1_carry ));
 XOR2_X2 \M2/stage3/gen_csa[1].FA0/HA1/_1_  (.A(\M2/sums2 [3]),
    .B(\M2/prodm3 [1]),
    .Z(\M2/stage3/gen_csa[1].FA0/ha1_sum ));
 AND2_X1 \M2/stage3/gen_csa[1].FA0/HA2/_0_  (.A1(\M2/stage3/gen_csa[1].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M2/stage3/gen_csa[1].FA0/ha2_carry ));
 XOR2_X1 \M2/stage3/gen_csa[1].FA0/HA2/_1_  (.A(\M2/stage3/gen_csa[1].FA0/ha1_sum ),
    .B(ground),
    .Z(\M2/stage3/sum0 [1]));
 OR2_X1 \M2/stage3/gen_csa[1].FA0/_0_  (.A1(\M2/stage3/gen_csa[1].FA0/ha1_carry ),
    .A2(\M2/stage3/gen_csa[1].FA0/ha2_carry ),
    .ZN(\M2/stage3/carry0 [1]));
 AND2_X1 \M2/stage3/gen_csa[1].FA1/HA1/_0_  (.A1(\M2/sums2 [3]),
    .A2(\M2/prodm3 [1]),
    .ZN(\M2/stage3/gen_csa[1].FA1/ha1_carry ));
 XOR2_X2 \M2/stage3/gen_csa[1].FA1/HA1/_1_  (.A(\M2/sums2 [3]),
    .B(\M2/prodm3 [1]),
    .Z(\M2/stage3/gen_csa[1].FA1/ha1_sum ));
 AND2_X1 \M2/stage3/gen_csa[1].FA1/HA2/_0_  (.A1(\M2/stage3/gen_csa[1].FA1/ha1_sum ),
    .A2(\M2/stage3/_03_ ),
    .ZN(\M2/stage3/gen_csa[1].FA1/ha2_carry ));
 XOR2_X1 \M2/stage3/gen_csa[1].FA1/HA2/_1_  (.A(\M2/stage3/gen_csa[1].FA1/ha1_sum ),
    .B(\M2/stage3/_03_ ),
    .Z(\M2/stage3/sum1 [1]));
 OR2_X1 \M2/stage3/gen_csa[1].FA1/_0_  (.A1(\M2/stage3/gen_csa[1].FA1/ha1_carry ),
    .A2(\M2/stage3/gen_csa[1].FA1/ha2_carry ),
    .ZN(\M2/stage3/carry1 [1]));
 AND2_X1 \M2/stage3/gen_csa[2].FA0/HA1/_0_  (.A1(\M2/cnet ),
    .A2(\M2/prodm3 [2]),
    .ZN(\M2/stage3/gen_csa[2].FA0/ha1_carry ));
 XOR2_X2 \M2/stage3/gen_csa[2].FA0/HA1/_1_  (.A(\M2/cnet ),
    .B(\M2/prodm3 [2]),
    .Z(\M2/stage3/gen_csa[2].FA0/ha1_sum ));
 AND2_X1 \M2/stage3/gen_csa[2].FA0/HA2/_0_  (.A1(\M2/stage3/gen_csa[2].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M2/stage3/gen_csa[2].FA0/ha2_carry ));
 XOR2_X1 \M2/stage3/gen_csa[2].FA0/HA2/_1_  (.A(\M2/stage3/gen_csa[2].FA0/ha1_sum ),
    .B(ground),
    .Z(\M2/stage3/sum0 [2]));
 OR2_X1 \M2/stage3/gen_csa[2].FA0/_0_  (.A1(\M2/stage3/gen_csa[2].FA0/ha1_carry ),
    .A2(\M2/stage3/gen_csa[2].FA0/ha2_carry ),
    .ZN(\M2/stage3/carry0 [2]));
 AND2_X1 \M2/stage3/gen_csa[2].FA1/HA1/_0_  (.A1(\M2/cnet ),
    .A2(\M2/prodm3 [2]),
    .ZN(\M2/stage3/gen_csa[2].FA1/ha1_carry ));
 XOR2_X2 \M2/stage3/gen_csa[2].FA1/HA1/_1_  (.A(\M2/cnet ),
    .B(\M2/prodm3 [2]),
    .Z(\M2/stage3/gen_csa[2].FA1/ha1_sum ));
 AND2_X1 \M2/stage3/gen_csa[2].FA1/HA2/_0_  (.A1(\M2/stage3/gen_csa[2].FA1/ha1_sum ),
    .A2(\M2/stage3/_03_ ),
    .ZN(\M2/stage3/gen_csa[2].FA1/ha2_carry ));
 XOR2_X1 \M2/stage3/gen_csa[2].FA1/HA2/_1_  (.A(\M2/stage3/gen_csa[2].FA1/ha1_sum ),
    .B(\M2/stage3/_03_ ),
    .Z(\M2/stage3/sum1 [2]));
 OR2_X1 \M2/stage3/gen_csa[2].FA1/_0_  (.A1(\M2/stage3/gen_csa[2].FA1/ha1_carry ),
    .A2(\M2/stage3/gen_csa[2].FA1/ha2_carry ),
    .ZN(\M2/stage3/carry1 [2]));
 AND2_X1 \M2/stage3/gen_csa[3].FA0/HA1/_0_  (.A1(ground),
    .A2(\M2/prodm3 [3]),
    .ZN(\M2/stage3/gen_csa[3].FA0/ha1_carry ));
 XOR2_X2 \M2/stage3/gen_csa[3].FA0/HA1/_1_  (.A(ground),
    .B(\M2/prodm3 [3]),
    .Z(\M2/stage3/gen_csa[3].FA0/ha1_sum ));
 AND2_X1 \M2/stage3/gen_csa[3].FA0/HA2/_0_  (.A1(\M2/stage3/gen_csa[3].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M2/stage3/gen_csa[3].FA0/ha2_carry ));
 XOR2_X1 \M2/stage3/gen_csa[3].FA0/HA2/_1_  (.A(\M2/stage3/gen_csa[3].FA0/ha1_sum ),
    .B(ground),
    .Z(\M2/stage3/sum0 [3]));
 OR2_X1 \M2/stage3/gen_csa[3].FA0/_0_  (.A1(\M2/stage3/gen_csa[3].FA0/ha1_carry ),
    .A2(\M2/stage3/gen_csa[3].FA0/ha2_carry ),
    .ZN(\M2/stage3/carry0 [3]));
 AND2_X1 \M2/stage3/gen_csa[3].FA1/HA1/_0_  (.A1(ground),
    .A2(\M2/prodm3 [3]),
    .ZN(\M2/stage3/gen_csa[3].FA1/ha1_carry ));
 XOR2_X2 \M2/stage3/gen_csa[3].FA1/HA1/_1_  (.A(ground),
    .B(\M2/prodm3 [3]),
    .Z(\M2/stage3/gen_csa[3].FA1/ha1_sum ));
 AND2_X1 \M2/stage3/gen_csa[3].FA1/HA2/_0_  (.A1(\M2/stage3/gen_csa[3].FA1/ha1_sum ),
    .A2(\M2/stage3/_03_ ),
    .ZN(\M2/stage3/gen_csa[3].FA1/ha2_carry ));
 XOR2_X1 \M2/stage3/gen_csa[3].FA1/HA2/_1_  (.A(\M2/stage3/gen_csa[3].FA1/ha1_sum ),
    .B(\M2/stage3/_03_ ),
    .Z(\M2/stage3/sum1 [3]));
 OR2_X1 \M2/stage3/gen_csa[3].FA1/_0_  (.A1(\M2/stage3/gen_csa[3].FA1/ha1_carry ),
    .A2(\M2/stage3/gen_csa[3].FA1/ha2_carry ),
    .ZN(\M2/stage3/carry1 [3]));
 AND2_X1 \M3/M0/HA0/_0_  (.A1(\M3/M0/a0b1 ),
    .A2(\M3/M0/a1b0 ),
    .ZN(\M3/M0/carry ));
 XOR2_X1 \M3/M0/HA0/_1_  (.A(\M3/M0/a0b1 ),
    .B(\M3/M0/a1b0 ),
    .Z(prodm3[1]));
 AND2_X1 \M3/M0/HA1/_0_  (.A1(\M3/M0/a1b1 ),
    .A2(\M3/M0/carry ),
    .ZN(\M3/prodm0 [3]));
 XOR2_X2 \M3/M0/HA1/_1_  (.A(\M3/M0/a1b1 ),
    .B(\M3/M0/carry ),
    .Z(\M3/prodm0 [2]));
 AND2_X1 \M3/M0/_0_  (.A1(a[5]),
    .A2(b[5]),
    .ZN(\M3/M0/a1b1 ));
 AND2_X1 \M3/M0/_1_  (.A1(b[5]),
    .A2(a[4]),
    .ZN(\M3/M0/a0b1 ));
 AND2_X1 \M3/M0/_2_  (.A1(a[5]),
    .A2(b[4]),
    .ZN(\M3/M0/a1b0 ));
 AND2_X1 \M3/M0/_3_  (.A1(a[4]),
    .A2(b[4]),
    .ZN(prodm3[0]));
 AND2_X1 \M3/M1/HA0/_0_  (.A1(\M3/M1/a0b1 ),
    .A2(\M3/M1/a1b0 ),
    .ZN(\M3/M1/carry ));
 XOR2_X2 \M3/M1/HA0/_1_  (.A(\M3/M1/a0b1 ),
    .B(\M3/M1/a1b0 ),
    .Z(\M3/prodm1 [1]));
 AND2_X1 \M3/M1/HA1/_0_  (.A1(\M3/M1/a1b1 ),
    .A2(\M3/M1/carry ),
    .ZN(\M3/prodm1 [3]));
 XOR2_X2 \M3/M1/HA1/_1_  (.A(\M3/M1/a1b1 ),
    .B(\M3/M1/carry ),
    .Z(\M3/prodm1 [2]));
 AND2_X1 \M3/M1/_0_  (.A1(a[5]),
    .A2(b[7]),
    .ZN(\M3/M1/a1b1 ));
 AND2_X1 \M3/M1/_1_  (.A1(b[7]),
    .A2(a[4]),
    .ZN(\M3/M1/a0b1 ));
 AND2_X1 \M3/M1/_2_  (.A1(a[5]),
    .A2(b[6]),
    .ZN(\M3/M1/a1b0 ));
 AND2_X1 \M3/M1/_3_  (.A1(a[4]),
    .A2(b[6]),
    .ZN(\M3/prodm1 [0]));
 AND2_X1 \M3/M2/HA0/_0_  (.A1(\M3/M2/a0b1 ),
    .A2(\M3/M2/a1b0 ),
    .ZN(\M3/M2/carry ));
 XOR2_X2 \M3/M2/HA0/_1_  (.A(\M3/M2/a0b1 ),
    .B(\M3/M2/a1b0 ),
    .Z(\M3/prodm2 [1]));
 AND2_X1 \M3/M2/HA1/_0_  (.A1(\M3/M2/a1b1 ),
    .A2(\M3/M2/carry ),
    .ZN(\M3/prodm2 [3]));
 XOR2_X2 \M3/M2/HA1/_1_  (.A(\M3/M2/a1b1 ),
    .B(\M3/M2/carry ),
    .Z(\M3/prodm2 [2]));
 AND2_X1 \M3/M2/_0_  (.A1(a[7]),
    .A2(b[5]),
    .ZN(\M3/M2/a1b1 ));
 AND2_X1 \M3/M2/_1_  (.A1(b[5]),
    .A2(a[6]),
    .ZN(\M3/M2/a0b1 ));
 AND2_X1 \M3/M2/_2_  (.A1(a[7]),
    .A2(b[4]),
    .ZN(\M3/M2/a1b0 ));
 AND2_X1 \M3/M2/_3_  (.A1(a[6]),
    .A2(b[4]),
    .ZN(\M3/prodm2 [0]));
 AND2_X1 \M3/M3/HA0/_0_  (.A1(\M3/M3/a0b1 ),
    .A2(\M3/M3/a1b0 ),
    .ZN(\M3/M3/carry ));
 XOR2_X2 \M3/M3/HA0/_1_  (.A(\M3/M3/a0b1 ),
    .B(\M3/M3/a1b0 ),
    .Z(\M3/prodm3 [1]));
 AND2_X1 \M3/M3/HA1/_0_  (.A1(\M3/M3/a1b1 ),
    .A2(\M3/M3/carry ),
    .ZN(\M3/prodm3 [3]));
 XOR2_X2 \M3/M3/HA1/_1_  (.A(\M3/M3/a1b1 ),
    .B(\M3/M3/carry ),
    .Z(\M3/prodm3 [2]));
 AND2_X1 \M3/M3/_0_  (.A1(a[7]),
    .A2(b[7]),
    .ZN(\M3/M3/a1b1 ));
 AND2_X1 \M3/M3/_1_  (.A1(b[7]),
    .A2(a[6]),
    .ZN(\M3/M3/a0b1 ));
 AND2_X1 \M3/M3/_2_  (.A1(a[7]),
    .A2(b[6]),
    .ZN(\M3/M3/a1b0 ));
 AND2_X1 \M3/M3/_3_  (.A1(a[6]),
    .A2(b[6]),
    .ZN(\M3/prodm3 [0]));
 OR2_X2 \M3/_0_  (.A1(\M3/c1 ),
    .A2(\M3/c2 ),
    .ZN(\M3/cnet ));
 AND2_X1 \M3/stage1/FA1_0/HA1/_0_  (.A1(\M3/prodm1 [0]),
    .A2(\M3/prodm2 [0]),
    .ZN(\M3/stage1/FA1_0/ha1_carry ));
 XOR2_X2 \M3/stage1/FA1_0/HA1/_1_  (.A(\M3/prodm1 [0]),
    .B(\M3/prodm2 [0]),
    .Z(\M3/stage1/FA1_0/ha1_sum ));
 AND2_X1 \M3/stage1/FA1_0/HA2/_0_  (.A1(\M3/stage1/FA1_0/ha1_sum ),
    .A2(\M3/stage1/_03_ ),
    .ZN(\M3/stage1/FA1_0/ha2_carry ));
 XOR2_X1 \M3/stage1/FA1_0/HA2/_1_  (.A(\M3/stage1/FA1_0/ha1_sum ),
    .B(\M3/stage1/_03_ ),
    .Z(\M3/stage1/sum1 [0]));
 OR2_X1 \M3/stage1/FA1_0/_0_  (.A1(\M3/stage1/FA1_0/ha1_carry ),
    .A2(\M3/stage1/FA1_0/ha2_carry ),
    .ZN(\M3/stage1/carry1 [0]));
 AND2_X1 \M3/stage1/HA0_0/_0_  (.A1(\M3/prodm1 [0]),
    .A2(\M3/prodm2 [0]),
    .ZN(\M3/stage1/carry0 [0]));
 XOR2_X1 \M3/stage1/HA0_0/_1_  (.A(\M3/prodm1 [0]),
    .B(\M3/prodm2 [0]),
    .Z(\M3/stage1/sum0 [0]));
 INV_X2 \M3/stage1/_04_  (.A(ground),
    .ZN(\M3/stage1/_03_ ));
 MUX2_X2 \M3/stage1/_05_  (.A(\M3/stage1/sum0 [0]),
    .B(\M3/stage1/sum1 [0]),
    .S(ground),
    .Z(\M3/sums1 [0]));
 MUX2_X1 \M3/stage1/_06_  (.A(\M3/stage1/carry0 [0]),
    .B(\M3/stage1/carry1 [0]),
    .S(ground),
    .Z(\M3/stage1/_00_ ));
 MUX2_X2 \M3/stage1/_07_  (.A(\M3/stage1/sum0 [1]),
    .B(\M3/stage1/sum1 [1]),
    .S(\M3/stage1/_00_ ),
    .Z(\M3/sums1 [1]));
 MUX2_X1 \M3/stage1/_08_  (.A(\M3/stage1/carry0 [1]),
    .B(\M3/stage1/carry1 [1]),
    .S(\M3/stage1/_00_ ),
    .Z(\M3/stage1/_01_ ));
 MUX2_X2 \M3/stage1/_09_  (.A(\M3/stage1/sum0 [2]),
    .B(\M3/stage1/sum1 [2]),
    .S(\M3/stage1/_01_ ),
    .Z(\M3/sums1 [2]));
 MUX2_X1 \M3/stage1/_10_  (.A(\M3/stage1/carry0 [2]),
    .B(\M3/stage1/carry1 [2]),
    .S(\M3/stage1/_01_ ),
    .Z(\M3/stage1/_02_ ));
 MUX2_X2 \M3/stage1/_11_  (.A(\M3/stage1/sum0 [3]),
    .B(\M3/stage1/sum1 [3]),
    .S(\M3/stage1/_02_ ),
    .Z(\M3/sums1 [3]));
 MUX2_X1 \M3/stage1/_12_  (.A(\M3/stage1/carry0 [3]),
    .B(\M3/stage1/carry1 [3]),
    .S(\M3/stage1/_02_ ),
    .Z(\M3/c1 ));
 AND2_X1 \M3/stage1/gen_csa[1].FA0/HA1/_0_  (.A1(\M3/prodm1 [1]),
    .A2(\M3/prodm2 [1]),
    .ZN(\M3/stage1/gen_csa[1].FA0/ha1_carry ));
 XOR2_X2 \M3/stage1/gen_csa[1].FA0/HA1/_1_  (.A(\M3/prodm1 [1]),
    .B(\M3/prodm2 [1]),
    .Z(\M3/stage1/gen_csa[1].FA0/ha1_sum ));
 AND2_X1 \M3/stage1/gen_csa[1].FA0/HA2/_0_  (.A1(\M3/stage1/gen_csa[1].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M3/stage1/gen_csa[1].FA0/ha2_carry ));
 XOR2_X1 \M3/stage1/gen_csa[1].FA0/HA2/_1_  (.A(\M3/stage1/gen_csa[1].FA0/ha1_sum ),
    .B(ground),
    .Z(\M3/stage1/sum0 [1]));
 OR2_X1 \M3/stage1/gen_csa[1].FA0/_0_  (.A1(\M3/stage1/gen_csa[1].FA0/ha1_carry ),
    .A2(\M3/stage1/gen_csa[1].FA0/ha2_carry ),
    .ZN(\M3/stage1/carry0 [1]));
 AND2_X1 \M3/stage1/gen_csa[1].FA1/HA1/_0_  (.A1(\M3/prodm1 [1]),
    .A2(\M3/prodm2 [1]),
    .ZN(\M3/stage1/gen_csa[1].FA1/ha1_carry ));
 XOR2_X2 \M3/stage1/gen_csa[1].FA1/HA1/_1_  (.A(\M3/prodm1 [1]),
    .B(\M3/prodm2 [1]),
    .Z(\M3/stage1/gen_csa[1].FA1/ha1_sum ));
 AND2_X1 \M3/stage1/gen_csa[1].FA1/HA2/_0_  (.A1(\M3/stage1/gen_csa[1].FA1/ha1_sum ),
    .A2(\M3/stage1/_03_ ),
    .ZN(\M3/stage1/gen_csa[1].FA1/ha2_carry ));
 XOR2_X1 \M3/stage1/gen_csa[1].FA1/HA2/_1_  (.A(\M3/stage1/gen_csa[1].FA1/ha1_sum ),
    .B(\M3/stage1/_03_ ),
    .Z(\M3/stage1/sum1 [1]));
 OR2_X1 \M3/stage1/gen_csa[1].FA1/_0_  (.A1(\M3/stage1/gen_csa[1].FA1/ha1_carry ),
    .A2(\M3/stage1/gen_csa[1].FA1/ha2_carry ),
    .ZN(\M3/stage1/carry1 [1]));
 AND2_X1 \M3/stage1/gen_csa[2].FA0/HA1/_0_  (.A1(\M3/prodm1 [2]),
    .A2(\M3/prodm2 [2]),
    .ZN(\M3/stage1/gen_csa[2].FA0/ha1_carry ));
 XOR2_X2 \M3/stage1/gen_csa[2].FA0/HA1/_1_  (.A(\M3/prodm1 [2]),
    .B(\M3/prodm2 [2]),
    .Z(\M3/stage1/gen_csa[2].FA0/ha1_sum ));
 AND2_X1 \M3/stage1/gen_csa[2].FA0/HA2/_0_  (.A1(\M3/stage1/gen_csa[2].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M3/stage1/gen_csa[2].FA0/ha2_carry ));
 XOR2_X1 \M3/stage1/gen_csa[2].FA0/HA2/_1_  (.A(\M3/stage1/gen_csa[2].FA0/ha1_sum ),
    .B(ground),
    .Z(\M3/stage1/sum0 [2]));
 OR2_X1 \M3/stage1/gen_csa[2].FA0/_0_  (.A1(\M3/stage1/gen_csa[2].FA0/ha1_carry ),
    .A2(\M3/stage1/gen_csa[2].FA0/ha2_carry ),
    .ZN(\M3/stage1/carry0 [2]));
 AND2_X1 \M3/stage1/gen_csa[2].FA1/HA1/_0_  (.A1(\M3/prodm1 [2]),
    .A2(\M3/prodm2 [2]),
    .ZN(\M3/stage1/gen_csa[2].FA1/ha1_carry ));
 XOR2_X2 \M3/stage1/gen_csa[2].FA1/HA1/_1_  (.A(\M3/prodm1 [2]),
    .B(\M3/prodm2 [2]),
    .Z(\M3/stage1/gen_csa[2].FA1/ha1_sum ));
 AND2_X1 \M3/stage1/gen_csa[2].FA1/HA2/_0_  (.A1(\M3/stage1/gen_csa[2].FA1/ha1_sum ),
    .A2(\M3/stage1/_03_ ),
    .ZN(\M3/stage1/gen_csa[2].FA1/ha2_carry ));
 XOR2_X1 \M3/stage1/gen_csa[2].FA1/HA2/_1_  (.A(\M3/stage1/gen_csa[2].FA1/ha1_sum ),
    .B(\M3/stage1/_03_ ),
    .Z(\M3/stage1/sum1 [2]));
 OR2_X1 \M3/stage1/gen_csa[2].FA1/_0_  (.A1(\M3/stage1/gen_csa[2].FA1/ha1_carry ),
    .A2(\M3/stage1/gen_csa[2].FA1/ha2_carry ),
    .ZN(\M3/stage1/carry1 [2]));
 AND2_X1 \M3/stage1/gen_csa[3].FA0/HA1/_0_  (.A1(\M3/prodm1 [3]),
    .A2(\M3/prodm2 [3]),
    .ZN(\M3/stage1/gen_csa[3].FA0/ha1_carry ));
 XOR2_X2 \M3/stage1/gen_csa[3].FA0/HA1/_1_  (.A(\M3/prodm1 [3]),
    .B(\M3/prodm2 [3]),
    .Z(\M3/stage1/gen_csa[3].FA0/ha1_sum ));
 AND2_X1 \M3/stage1/gen_csa[3].FA0/HA2/_0_  (.A1(\M3/stage1/gen_csa[3].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M3/stage1/gen_csa[3].FA0/ha2_carry ));
 XOR2_X1 \M3/stage1/gen_csa[3].FA0/HA2/_1_  (.A(\M3/stage1/gen_csa[3].FA0/ha1_sum ),
    .B(ground),
    .Z(\M3/stage1/sum0 [3]));
 OR2_X1 \M3/stage1/gen_csa[3].FA0/_0_  (.A1(\M3/stage1/gen_csa[3].FA0/ha1_carry ),
    .A2(\M3/stage1/gen_csa[3].FA0/ha2_carry ),
    .ZN(\M3/stage1/carry0 [3]));
 AND2_X1 \M3/stage1/gen_csa[3].FA1/HA1/_0_  (.A1(\M3/prodm1 [3]),
    .A2(\M3/prodm2 [3]),
    .ZN(\M3/stage1/gen_csa[3].FA1/ha1_carry ));
 XOR2_X2 \M3/stage1/gen_csa[3].FA1/HA1/_1_  (.A(\M3/prodm1 [3]),
    .B(\M3/prodm2 [3]),
    .Z(\M3/stage1/gen_csa[3].FA1/ha1_sum ));
 AND2_X1 \M3/stage1/gen_csa[3].FA1/HA2/_0_  (.A1(\M3/stage1/gen_csa[3].FA1/ha1_sum ),
    .A2(\M3/stage1/_03_ ),
    .ZN(\M3/stage1/gen_csa[3].FA1/ha2_carry ));
 XOR2_X1 \M3/stage1/gen_csa[3].FA1/HA2/_1_  (.A(\M3/stage1/gen_csa[3].FA1/ha1_sum ),
    .B(\M3/stage1/_03_ ),
    .Z(\M3/stage1/sum1 [3]));
 OR2_X1 \M3/stage1/gen_csa[3].FA1/_0_  (.A1(\M3/stage1/gen_csa[3].FA1/ha1_carry ),
    .A2(\M3/stage1/gen_csa[3].FA1/ha2_carry ),
    .ZN(\M3/stage1/carry1 [3]));
 AND2_X1 \M3/stage2/FA1_0/HA1/_0_  (.A1(\M3/prodm0 [2]),
    .A2(\M3/sums1 [0]),
    .ZN(\M3/stage2/FA1_0/ha1_carry ));
 XOR2_X2 \M3/stage2/FA1_0/HA1/_1_  (.A(\M3/prodm0 [2]),
    .B(\M3/sums1 [0]),
    .Z(\M3/stage2/FA1_0/ha1_sum ));
 AND2_X1 \M3/stage2/FA1_0/HA2/_0_  (.A1(\M3/stage2/FA1_0/ha1_sum ),
    .A2(\M3/stage2/_03_ ),
    .ZN(\M3/stage2/FA1_0/ha2_carry ));
 XOR2_X1 \M3/stage2/FA1_0/HA2/_1_  (.A(\M3/stage2/FA1_0/ha1_sum ),
    .B(\M3/stage2/_03_ ),
    .Z(\M3/stage2/sum1 [0]));
 OR2_X1 \M3/stage2/FA1_0/_0_  (.A1(\M3/stage2/FA1_0/ha1_carry ),
    .A2(\M3/stage2/FA1_0/ha2_carry ),
    .ZN(\M3/stage2/carry1 [0]));
 AND2_X1 \M3/stage2/HA0_0/_0_  (.A1(\M3/prodm0 [2]),
    .A2(\M3/sums1 [0]),
    .ZN(\M3/stage2/carry0 [0]));
 XOR2_X1 \M3/stage2/HA0_0/_1_  (.A(\M3/prodm0 [2]),
    .B(\M3/sums1 [0]),
    .Z(\M3/stage2/sum0 [0]));
 INV_X2 \M3/stage2/_04_  (.A(ground),
    .ZN(\M3/stage2/_03_ ));
 MUX2_X1 \M3/stage2/_05_  (.A(\M3/stage2/sum0 [0]),
    .B(\M3/stage2/sum1 [0]),
    .S(ground),
    .Z(prodm3[2]));
 MUX2_X1 \M3/stage2/_06_  (.A(\M3/stage2/carry0 [0]),
    .B(\M3/stage2/carry1 [0]),
    .S(ground),
    .Z(\M3/stage2/_00_ ));
 MUX2_X1 \M3/stage2/_07_  (.A(\M3/stage2/sum0 [1]),
    .B(\M3/stage2/sum1 [1]),
    .S(\M3/stage2/_00_ ),
    .Z(prodm3[3]));
 MUX2_X1 \M3/stage2/_08_  (.A(\M3/stage2/carry0 [1]),
    .B(\M3/stage2/carry1 [1]),
    .S(\M3/stage2/_00_ ),
    .Z(\M3/stage2/_01_ ));
 MUX2_X1 \M3/stage2/_09_  (.A(\M3/stage2/sum0 [2]),
    .B(\M3/stage2/sum1 [2]),
    .S(\M3/stage2/_01_ ),
    .Z(\M3/sums2 [2]));
 MUX2_X1 \M3/stage2/_10_  (.A(\M3/stage2/carry0 [2]),
    .B(\M3/stage2/carry1 [2]),
    .S(\M3/stage2/_01_ ),
    .Z(\M3/stage2/_02_ ));
 MUX2_X2 \M3/stage2/_11_  (.A(\M3/stage2/sum0 [3]),
    .B(\M3/stage2/sum1 [3]),
    .S(\M3/stage2/_02_ ),
    .Z(\M3/sums2 [3]));
 MUX2_X1 \M3/stage2/_12_  (.A(\M3/stage2/carry0 [3]),
    .B(\M3/stage2/carry1 [3]),
    .S(\M3/stage2/_02_ ),
    .Z(\M3/c2 ));
 AND2_X1 \M3/stage2/gen_csa[1].FA0/HA1/_0_  (.A1(\M3/prodm0 [3]),
    .A2(\M3/sums1 [1]),
    .ZN(\M3/stage2/gen_csa[1].FA0/ha1_carry ));
 XOR2_X2 \M3/stage2/gen_csa[1].FA0/HA1/_1_  (.A(\M3/prodm0 [3]),
    .B(\M3/sums1 [1]),
    .Z(\M3/stage2/gen_csa[1].FA0/ha1_sum ));
 AND2_X1 \M3/stage2/gen_csa[1].FA0/HA2/_0_  (.A1(\M3/stage2/gen_csa[1].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M3/stage2/gen_csa[1].FA0/ha2_carry ));
 XOR2_X1 \M3/stage2/gen_csa[1].FA0/HA2/_1_  (.A(\M3/stage2/gen_csa[1].FA0/ha1_sum ),
    .B(ground),
    .Z(\M3/stage2/sum0 [1]));
 OR2_X1 \M3/stage2/gen_csa[1].FA0/_0_  (.A1(\M3/stage2/gen_csa[1].FA0/ha1_carry ),
    .A2(\M3/stage2/gen_csa[1].FA0/ha2_carry ),
    .ZN(\M3/stage2/carry0 [1]));
 AND2_X1 \M3/stage2/gen_csa[1].FA1/HA1/_0_  (.A1(\M3/prodm0 [3]),
    .A2(\M3/sums1 [1]),
    .ZN(\M3/stage2/gen_csa[1].FA1/ha1_carry ));
 XOR2_X2 \M3/stage2/gen_csa[1].FA1/HA1/_1_  (.A(\M3/prodm0 [3]),
    .B(\M3/sums1 [1]),
    .Z(\M3/stage2/gen_csa[1].FA1/ha1_sum ));
 AND2_X1 \M3/stage2/gen_csa[1].FA1/HA2/_0_  (.A1(\M3/stage2/gen_csa[1].FA1/ha1_sum ),
    .A2(\M3/stage2/_03_ ),
    .ZN(\M3/stage2/gen_csa[1].FA1/ha2_carry ));
 XOR2_X1 \M3/stage2/gen_csa[1].FA1/HA2/_1_  (.A(\M3/stage2/gen_csa[1].FA1/ha1_sum ),
    .B(\M3/stage2/_03_ ),
    .Z(\M3/stage2/sum1 [1]));
 OR2_X1 \M3/stage2/gen_csa[1].FA1/_0_  (.A1(\M3/stage2/gen_csa[1].FA1/ha1_carry ),
    .A2(\M3/stage2/gen_csa[1].FA1/ha2_carry ),
    .ZN(\M3/stage2/carry1 [1]));
 AND2_X1 \M3/stage2/gen_csa[2].FA0/HA1/_0_  (.A1(ground),
    .A2(\M3/sums1 [2]),
    .ZN(\M3/stage2/gen_csa[2].FA0/ha1_carry ));
 XOR2_X2 \M3/stage2/gen_csa[2].FA0/HA1/_1_  (.A(ground),
    .B(\M3/sums1 [2]),
    .Z(\M3/stage2/gen_csa[2].FA0/ha1_sum ));
 AND2_X1 \M3/stage2/gen_csa[2].FA0/HA2/_0_  (.A1(\M3/stage2/gen_csa[2].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M3/stage2/gen_csa[2].FA0/ha2_carry ));
 XOR2_X1 \M3/stage2/gen_csa[2].FA0/HA2/_1_  (.A(\M3/stage2/gen_csa[2].FA0/ha1_sum ),
    .B(ground),
    .Z(\M3/stage2/sum0 [2]));
 OR2_X1 \M3/stage2/gen_csa[2].FA0/_0_  (.A1(\M3/stage2/gen_csa[2].FA0/ha1_carry ),
    .A2(\M3/stage2/gen_csa[2].FA0/ha2_carry ),
    .ZN(\M3/stage2/carry0 [2]));
 AND2_X1 \M3/stage2/gen_csa[2].FA1/HA1/_0_  (.A1(ground),
    .A2(\M3/sums1 [2]),
    .ZN(\M3/stage2/gen_csa[2].FA1/ha1_carry ));
 XOR2_X2 \M3/stage2/gen_csa[2].FA1/HA1/_1_  (.A(ground),
    .B(\M3/sums1 [2]),
    .Z(\M3/stage2/gen_csa[2].FA1/ha1_sum ));
 AND2_X1 \M3/stage2/gen_csa[2].FA1/HA2/_0_  (.A1(\M3/stage2/gen_csa[2].FA1/ha1_sum ),
    .A2(\M3/stage2/_03_ ),
    .ZN(\M3/stage2/gen_csa[2].FA1/ha2_carry ));
 XOR2_X1 \M3/stage2/gen_csa[2].FA1/HA2/_1_  (.A(\M3/stage2/gen_csa[2].FA1/ha1_sum ),
    .B(\M3/stage2/_03_ ),
    .Z(\M3/stage2/sum1 [2]));
 OR2_X1 \M3/stage2/gen_csa[2].FA1/_0_  (.A1(\M3/stage2/gen_csa[2].FA1/ha1_carry ),
    .A2(\M3/stage2/gen_csa[2].FA1/ha2_carry ),
    .ZN(\M3/stage2/carry1 [2]));
 AND2_X1 \M3/stage2/gen_csa[3].FA0/HA1/_0_  (.A1(ground),
    .A2(\M3/sums1 [3]),
    .ZN(\M3/stage2/gen_csa[3].FA0/ha1_carry ));
 XOR2_X2 \M3/stage2/gen_csa[3].FA0/HA1/_1_  (.A(ground),
    .B(\M3/sums1 [3]),
    .Z(\M3/stage2/gen_csa[3].FA0/ha1_sum ));
 AND2_X1 \M3/stage2/gen_csa[3].FA0/HA2/_0_  (.A1(\M3/stage2/gen_csa[3].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M3/stage2/gen_csa[3].FA0/ha2_carry ));
 XOR2_X1 \M3/stage2/gen_csa[3].FA0/HA2/_1_  (.A(\M3/stage2/gen_csa[3].FA0/ha1_sum ),
    .B(ground),
    .Z(\M3/stage2/sum0 [3]));
 OR2_X1 \M3/stage2/gen_csa[3].FA0/_0_  (.A1(\M3/stage2/gen_csa[3].FA0/ha1_carry ),
    .A2(\M3/stage2/gen_csa[3].FA0/ha2_carry ),
    .ZN(\M3/stage2/carry0 [3]));
 AND2_X1 \M3/stage2/gen_csa[3].FA1/HA1/_0_  (.A1(ground),
    .A2(\M3/sums1 [3]),
    .ZN(\M3/stage2/gen_csa[3].FA1/ha1_carry ));
 XOR2_X1 \M3/stage2/gen_csa[3].FA1/HA1/_1_  (.A(ground),
    .B(\M3/sums1 [3]),
    .Z(\M3/stage2/gen_csa[3].FA1/ha1_sum ));
 AND2_X1 \M3/stage2/gen_csa[3].FA1/HA2/_0_  (.A1(\M3/stage2/gen_csa[3].FA1/ha1_sum ),
    .A2(\M3/stage2/_03_ ),
    .ZN(\M3/stage2/gen_csa[3].FA1/ha2_carry ));
 XOR2_X1 \M3/stage2/gen_csa[3].FA1/HA2/_1_  (.A(\M3/stage2/gen_csa[3].FA1/ha1_sum ),
    .B(\M3/stage2/_03_ ),
    .Z(\M3/stage2/sum1 [3]));
 OR2_X1 \M3/stage2/gen_csa[3].FA1/_0_  (.A1(\M3/stage2/gen_csa[3].FA1/ha1_carry ),
    .A2(\M3/stage2/gen_csa[3].FA1/ha2_carry ),
    .ZN(\M3/stage2/carry1 [3]));
 AND2_X1 \M3/stage3/FA1_0/HA1/_0_  (.A1(\M3/sums2 [2]),
    .A2(\M3/prodm3 [0]),
    .ZN(\M3/stage3/FA1_0/ha1_carry ));
 XOR2_X1 \M3/stage3/FA1_0/HA1/_1_  (.A(\M3/sums2 [2]),
    .B(\M3/prodm3 [0]),
    .Z(\M3/stage3/FA1_0/ha1_sum ));
 AND2_X1 \M3/stage3/FA1_0/HA2/_0_  (.A1(\M3/stage3/FA1_0/ha1_sum ),
    .A2(\M3/stage3/_03_ ),
    .ZN(\M3/stage3/FA1_0/ha2_carry ));
 XOR2_X1 \M3/stage3/FA1_0/HA2/_1_  (.A(\M3/stage3/FA1_0/ha1_sum ),
    .B(\M3/stage3/_03_ ),
    .Z(\M3/stage3/sum1 [0]));
 OR2_X1 \M3/stage3/FA1_0/_0_  (.A1(\M3/stage3/FA1_0/ha1_carry ),
    .A2(\M3/stage3/FA1_0/ha2_carry ),
    .ZN(\M3/stage3/carry1 [0]));
 AND2_X1 \M3/stage3/HA0_0/_0_  (.A1(\M3/sums2 [2]),
    .A2(\M3/prodm3 [0]),
    .ZN(\M3/stage3/carry0 [0]));
 XOR2_X1 \M3/stage3/HA0_0/_1_  (.A(\M3/sums2 [2]),
    .B(\M3/prodm3 [0]),
    .Z(\M3/stage3/sum0 [0]));
 INV_X2 \M3/stage3/_04_  (.A(ground),
    .ZN(\M3/stage3/_03_ ));
 MUX2_X1 \M3/stage3/_05_  (.A(\M3/stage3/sum0 [0]),
    .B(\M3/stage3/sum1 [0]),
    .S(ground),
    .Z(prodm3[4]));
 MUX2_X1 \M3/stage3/_06_  (.A(\M3/stage3/carry0 [0]),
    .B(\M3/stage3/carry1 [0]),
    .S(ground),
    .Z(\M3/stage3/_00_ ));
 MUX2_X1 \M3/stage3/_07_  (.A(\M3/stage3/sum0 [1]),
    .B(\M3/stage3/sum1 [1]),
    .S(\M3/stage3/_00_ ),
    .Z(prodm3[5]));
 MUX2_X1 \M3/stage3/_08_  (.A(\M3/stage3/carry0 [1]),
    .B(\M3/stage3/carry1 [1]),
    .S(\M3/stage3/_00_ ),
    .Z(\M3/stage3/_01_ ));
 MUX2_X1 \M3/stage3/_09_  (.A(\M3/stage3/sum0 [2]),
    .B(\M3/stage3/sum1 [2]),
    .S(\M3/stage3/_01_ ),
    .Z(prodm3[6]));
 MUX2_X1 \M3/stage3/_10_  (.A(\M3/stage3/carry0 [2]),
    .B(\M3/stage3/carry1 [2]),
    .S(\M3/stage3/_01_ ),
    .Z(\M3/stage3/_02_ ));
 MUX2_X1 \M3/stage3/_11_  (.A(\M3/stage3/sum0 [3]),
    .B(\M3/stage3/sum1 [3]),
    .S(\M3/stage3/_02_ ),
    .Z(prodm3[7]));
 MUX2_X1 \M3/stage3/_12_  (.A(\M3/stage3/carry0 [3]),
    .B(\M3/stage3/carry1 [3]),
    .S(\M3/stage3/_02_ ),
    .Z(ov4));
 AND2_X1 \M3/stage3/gen_csa[1].FA0/HA1/_0_  (.A1(\M3/sums2 [3]),
    .A2(\M3/prodm3 [1]),
    .ZN(\M3/stage3/gen_csa[1].FA0/ha1_carry ));
 XOR2_X2 \M3/stage3/gen_csa[1].FA0/HA1/_1_  (.A(\M3/sums2 [3]),
    .B(\M3/prodm3 [1]),
    .Z(\M3/stage3/gen_csa[1].FA0/ha1_sum ));
 AND2_X1 \M3/stage3/gen_csa[1].FA0/HA2/_0_  (.A1(\M3/stage3/gen_csa[1].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M3/stage3/gen_csa[1].FA0/ha2_carry ));
 XOR2_X1 \M3/stage3/gen_csa[1].FA0/HA2/_1_  (.A(\M3/stage3/gen_csa[1].FA0/ha1_sum ),
    .B(ground),
    .Z(\M3/stage3/sum0 [1]));
 OR2_X1 \M3/stage3/gen_csa[1].FA0/_0_  (.A1(\M3/stage3/gen_csa[1].FA0/ha1_carry ),
    .A2(\M3/stage3/gen_csa[1].FA0/ha2_carry ),
    .ZN(\M3/stage3/carry0 [1]));
 AND2_X1 \M3/stage3/gen_csa[1].FA1/HA1/_0_  (.A1(\M3/sums2 [3]),
    .A2(\M3/prodm3 [1]),
    .ZN(\M3/stage3/gen_csa[1].FA1/ha1_carry ));
 XOR2_X2 \M3/stage3/gen_csa[1].FA1/HA1/_1_  (.A(\M3/sums2 [3]),
    .B(\M3/prodm3 [1]),
    .Z(\M3/stage3/gen_csa[1].FA1/ha1_sum ));
 AND2_X1 \M3/stage3/gen_csa[1].FA1/HA2/_0_  (.A1(\M3/stage3/gen_csa[1].FA1/ha1_sum ),
    .A2(\M3/stage3/_03_ ),
    .ZN(\M3/stage3/gen_csa[1].FA1/ha2_carry ));
 XOR2_X1 \M3/stage3/gen_csa[1].FA1/HA2/_1_  (.A(\M3/stage3/gen_csa[1].FA1/ha1_sum ),
    .B(\M3/stage3/_03_ ),
    .Z(\M3/stage3/sum1 [1]));
 OR2_X1 \M3/stage3/gen_csa[1].FA1/_0_  (.A1(\M3/stage3/gen_csa[1].FA1/ha1_carry ),
    .A2(\M3/stage3/gen_csa[1].FA1/ha2_carry ),
    .ZN(\M3/stage3/carry1 [1]));
 AND2_X1 \M3/stage3/gen_csa[2].FA0/HA1/_0_  (.A1(\M3/cnet ),
    .A2(\M3/prodm3 [2]),
    .ZN(\M3/stage3/gen_csa[2].FA0/ha1_carry ));
 XOR2_X2 \M3/stage3/gen_csa[2].FA0/HA1/_1_  (.A(\M3/cnet ),
    .B(\M3/prodm3 [2]),
    .Z(\M3/stage3/gen_csa[2].FA0/ha1_sum ));
 AND2_X1 \M3/stage3/gen_csa[2].FA0/HA2/_0_  (.A1(\M3/stage3/gen_csa[2].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M3/stage3/gen_csa[2].FA0/ha2_carry ));
 XOR2_X1 \M3/stage3/gen_csa[2].FA0/HA2/_1_  (.A(\M3/stage3/gen_csa[2].FA0/ha1_sum ),
    .B(ground),
    .Z(\M3/stage3/sum0 [2]));
 OR2_X1 \M3/stage3/gen_csa[2].FA0/_0_  (.A1(\M3/stage3/gen_csa[2].FA0/ha1_carry ),
    .A2(\M3/stage3/gen_csa[2].FA0/ha2_carry ),
    .ZN(\M3/stage3/carry0 [2]));
 AND2_X1 \M3/stage3/gen_csa[2].FA1/HA1/_0_  (.A1(\M3/cnet ),
    .A2(\M3/prodm3 [2]),
    .ZN(\M3/stage3/gen_csa[2].FA1/ha1_carry ));
 XOR2_X2 \M3/stage3/gen_csa[2].FA1/HA1/_1_  (.A(\M3/cnet ),
    .B(\M3/prodm3 [2]),
    .Z(\M3/stage3/gen_csa[2].FA1/ha1_sum ));
 AND2_X1 \M3/stage3/gen_csa[2].FA1/HA2/_0_  (.A1(\M3/stage3/gen_csa[2].FA1/ha1_sum ),
    .A2(\M3/stage3/_03_ ),
    .ZN(\M3/stage3/gen_csa[2].FA1/ha2_carry ));
 XOR2_X1 \M3/stage3/gen_csa[2].FA1/HA2/_1_  (.A(\M3/stage3/gen_csa[2].FA1/ha1_sum ),
    .B(\M3/stage3/_03_ ),
    .Z(\M3/stage3/sum1 [2]));
 OR2_X1 \M3/stage3/gen_csa[2].FA1/_0_  (.A1(\M3/stage3/gen_csa[2].FA1/ha1_carry ),
    .A2(\M3/stage3/gen_csa[2].FA1/ha2_carry ),
    .ZN(\M3/stage3/carry1 [2]));
 AND2_X1 \M3/stage3/gen_csa[3].FA0/HA1/_0_  (.A1(ground),
    .A2(\M3/prodm3 [3]),
    .ZN(\M3/stage3/gen_csa[3].FA0/ha1_carry ));
 XOR2_X1 \M3/stage3/gen_csa[3].FA0/HA1/_1_  (.A(ground),
    .B(\M3/prodm3 [3]),
    .Z(\M3/stage3/gen_csa[3].FA0/ha1_sum ));
 AND2_X1 \M3/stage3/gen_csa[3].FA0/HA2/_0_  (.A1(\M3/stage3/gen_csa[3].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\M3/stage3/gen_csa[3].FA0/ha2_carry ));
 XOR2_X1 \M3/stage3/gen_csa[3].FA0/HA2/_1_  (.A(\M3/stage3/gen_csa[3].FA0/ha1_sum ),
    .B(ground),
    .Z(\M3/stage3/sum0 [3]));
 OR2_X1 \M3/stage3/gen_csa[3].FA0/_0_  (.A1(\M3/stage3/gen_csa[3].FA0/ha1_carry ),
    .A2(\M3/stage3/gen_csa[3].FA0/ha2_carry ),
    .ZN(\M3/stage3/carry0 [3]));
 AND2_X1 \M3/stage3/gen_csa[3].FA1/HA1/_0_  (.A1(ground),
    .A2(\M3/prodm3 [3]),
    .ZN(\M3/stage3/gen_csa[3].FA1/ha1_carry ));
 XOR2_X2 \M3/stage3/gen_csa[3].FA1/HA1/_1_  (.A(ground),
    .B(\M3/prodm3 [3]),
    .Z(\M3/stage3/gen_csa[3].FA1/ha1_sum ));
 AND2_X1 \M3/stage3/gen_csa[3].FA1/HA2/_0_  (.A1(\M3/stage3/gen_csa[3].FA1/ha1_sum ),
    .A2(\M3/stage3/_03_ ),
    .ZN(\M3/stage3/gen_csa[3].FA1/ha2_carry ));
 XOR2_X1 \M3/stage3/gen_csa[3].FA1/HA2/_1_  (.A(\M3/stage3/gen_csa[3].FA1/ha1_sum ),
    .B(\M3/stage3/_03_ ),
    .Z(\M3/stage3/sum1 [3]));
 OR2_X1 \M3/stage3/gen_csa[3].FA1/_0_  (.A1(\M3/stage3/gen_csa[3].FA1/ha1_carry ),
    .A2(\M3/stage3/gen_csa[3].FA1/ha2_carry ),
    .ZN(\M3/stage3/carry1 [3]));
 OR2_X2 _100_ (.A1(c1_s2),
    .A2(c2_s2),
    .ZN(_000_));
 DFF_X1 _101_ (.D(sums2[0]),
    .CK(clknet_3_5__leaf_clk),
    .Q(sum_s2[0]),
    .QN(_086_));
 DFF_X1 _102_ (.D(sums2[1]),
    .CK(clknet_3_5__leaf_clk),
    .Q(sum_s2[1]),
    .QN(_085_));
 DFF_X1 _103_ (.D(sums2[2]),
    .CK(clknet_3_2__leaf_clk),
    .Q(sum_s2[2]),
    .QN(_084_));
 DFF_X1 _104_ (.D(sums2[3]),
    .CK(clknet_3_4__leaf_clk),
    .Q(sum_s2[3]),
    .QN(_083_));
 DFF_X2 _105_ (.D(sums2[4]),
    .CK(clknet_3_4__leaf_clk),
    .Q(sum_s2[4]),
    .QN(_082_));
 DFF_X2 _106_ (.D(sums2[5]),
    .CK(clknet_3_6__leaf_clk),
    .Q(sum_s2[5]),
    .QN(_081_));
 DFF_X2 _107_ (.D(sums2[6]),
    .CK(clknet_3_3__leaf_clk),
    .Q(sum_s2[6]),
    .QN(_080_));
 DFF_X2 _108_ (.D(sums2[7]),
    .CK(clknet_3_3__leaf_clk),
    .Q(sum_s2[7]),
    .QN(_090_));
 DFF_X1 _109_ (.D(c1_s1),
    .CK(clknet_3_3__leaf_clk),
    .Q(c1_s2),
    .QN(_089_));
 DFF_X1 _110_ (.D(c2),
    .CK(clknet_3_3__leaf_clk),
    .Q(c2_s2),
    .QN(_088_));
 DFF_X1 _111_ (.D(prodm0_s2[0]),
    .CK(clknet_3_2__leaf_clk),
    .Q(prod[0]),
    .QN(_079_));
 DFF_X1 _112_ (.D(prodm0_s2[1]),
    .CK(clknet_3_0__leaf_clk),
    .Q(prod[1]),
    .QN(_078_));
 DFF_X1 _113_ (.D(prodm0_s2[2]),
    .CK(clknet_3_7__leaf_clk),
    .Q(prod[2]),
    .QN(_077_));
 DFF_X1 _114_ (.D(prodm0_s2[3]),
    .CK(clknet_3_7__leaf_clk),
    .Q(prod[3]),
    .QN(_076_));
 DFF_X1 _115_ (.D(sum_s2[0]),
    .CK(clknet_3_5__leaf_clk),
    .Q(prod[4]),
    .QN(_075_));
 DFF_X1 _116_ (.D(sum_s2[1]),
    .CK(clknet_3_5__leaf_clk),
    .Q(prod[5]),
    .QN(_074_));
 DFF_X1 _117_ (.D(sum_s2[2]),
    .CK(clknet_3_2__leaf_clk),
    .Q(prod[6]),
    .QN(_073_));
 DFF_X1 _118_ (.D(sum_s2[3]),
    .CK(clknet_3_1__leaf_clk),
    .Q(prod[7]),
    .QN(_072_));
 DFF_X1 _119_ (.D(sums3[0]),
    .CK(clknet_3_5__leaf_clk),
    .Q(prod[8]),
    .QN(_071_));
 DFF_X1 _120_ (.D(sums3[1]),
    .CK(clknet_3_6__leaf_clk),
    .Q(prod[9]),
    .QN(_070_));
 DFF_X1 _121_ (.D(sums3[2]),
    .CK(clknet_3_6__leaf_clk),
    .Q(prod[10]),
    .QN(_069_));
 DFF_X1 _122_ (.D(sums3[3]),
    .CK(clknet_3_2__leaf_clk),
    .Q(prod[11]),
    .QN(_068_));
 DFF_X1 _123_ (.D(sums3[4]),
    .CK(clknet_3_0__leaf_clk),
    .Q(prod[12]),
    .QN(_067_));
 DFF_X1 _124_ (.D(sums3[5]),
    .CK(clknet_3_0__leaf_clk),
    .Q(prod[13]),
    .QN(_066_));
 DFF_X1 _125_ (.D(sums3[6]),
    .CK(clknet_3_0__leaf_clk),
    .Q(prod[14]),
    .QN(_065_));
 DFF_X1 _126_ (.D(sums3[7]),
    .CK(clknet_3_2__leaf_clk),
    .Q(prod[15]),
    .QN(_087_));
 DFF_X1 _127_ (.D(prodm0_s1[0]),
    .CK(clknet_3_2__leaf_clk),
    .Q(prodm0_s2[0]),
    .QN(_064_));
 DFF_X1 _128_ (.D(prodm0_s1[1]),
    .CK(clknet_3_0__leaf_clk),
    .Q(prodm0_s2[1]),
    .QN(_063_));
 DFF_X1 _129_ (.D(prodm0_s1[2]),
    .CK(clknet_3_7__leaf_clk),
    .Q(prodm0_s2[2]),
    .QN(_062_));
 DFF_X1 _130_ (.D(prodm0_s1[3]),
    .CK(clknet_3_7__leaf_clk),
    .Q(prodm0_s2[3]),
    .QN(_061_));
 DFF_X1 _131_ (.D(prodm0_s1[4]),
    .CK(clknet_3_5__leaf_clk),
    .Q(prodm0_s2[4]),
    .QN(_060_));
 DFF_X1 _132_ (.D(prodm0_s1[5]),
    .CK(clknet_3_5__leaf_clk),
    .Q(prodm0_s2[5]),
    .QN(_059_));
 DFF_X1 _133_ (.D(prodm0_s1[6]),
    .CK(clknet_3_5__leaf_clk),
    .Q(prodm0_s2[6]),
    .QN(_058_));
 DFF_X1 _134_ (.D(prodm0_s1[7]),
    .CK(clknet_3_6__leaf_clk),
    .Q(prodm0_s2[7]),
    .QN(_091_));
 DFF_X2 _135_ (.D(prodm3_s1[0]),
    .CK(clknet_3_4__leaf_clk),
    .Q(prodm3_s2[0]),
    .QN(_057_));
 DFF_X2 _136_ (.D(prodm3_s1[1]),
    .CK(clknet_3_6__leaf_clk),
    .Q(prodm3_s2[1]),
    .QN(_056_));
 DFF_X2 _137_ (.D(prodm3_s1[2]),
    .CK(clknet_3_3__leaf_clk),
    .Q(prodm3_s2[2]),
    .QN(_055_));
 DFF_X2 _138_ (.D(prodm3_s1[3]),
    .CK(clknet_3_1__leaf_clk),
    .Q(prodm3_s2[3]),
    .QN(_054_));
 DFF_X2 _139_ (.D(prodm3_s1[4]),
    .CK(clknet_3_0__leaf_clk),
    .Q(prodm3_s2[4]),
    .QN(_053_));
 DFF_X2 _140_ (.D(prodm3_s1[5]),
    .CK(clknet_3_0__leaf_clk),
    .Q(prodm3_s2[5]),
    .QN(_052_));
 DFF_X2 _141_ (.D(prodm3_s1[6]),
    .CK(clknet_3_0__leaf_clk),
    .Q(prodm3_s2[6]),
    .QN(_051_));
 DFF_X2 _142_ (.D(prodm3_s1[7]),
    .CK(clknet_3_0__leaf_clk),
    .Q(prodm3_s2[7]),
    .QN(_092_));
 DFF_X1 _143_ (.D(c1),
    .CK(clknet_3_1__leaf_clk),
    .Q(c1_s1),
    .QN(_093_));
 DFF_X1 _144_ (.D(prodm0_s0[0]),
    .CK(clknet_3_6__leaf_clk),
    .Q(prodm0_s1[0]),
    .QN(_050_));
 DFF_X1 _145_ (.D(prodm0_s0[1]),
    .CK(clknet_3_0__leaf_clk),
    .Q(prodm0_s1[1]),
    .QN(_049_));
 DFF_X1 _146_ (.D(prodm0_s0[2]),
    .CK(clknet_3_7__leaf_clk),
    .Q(prodm0_s1[2]),
    .QN(_048_));
 DFF_X1 _147_ (.D(prodm0_s0[3]),
    .CK(clknet_3_7__leaf_clk),
    .Q(prodm0_s1[3]),
    .QN(_047_));
 DFF_X2 _148_ (.D(prodm0_s0[4]),
    .CK(clknet_3_5__leaf_clk),
    .Q(prodm0_s1[4]),
    .QN(_046_));
 DFF_X2 _149_ (.D(prodm0_s0[5]),
    .CK(clknet_3_5__leaf_clk),
    .Q(prodm0_s1[5]),
    .QN(_045_));
 DFF_X2 _150_ (.D(prodm0_s0[6]),
    .CK(clknet_3_5__leaf_clk),
    .Q(prodm0_s1[6]),
    .QN(_044_));
 DFF_X2 _151_ (.D(prodm0_s0[7]),
    .CK(clknet_3_6__leaf_clk),
    .Q(prodm0_s1[7]),
    .QN(_094_));
 DFF_X1 _152_ (.D(prodm3_s0[0]),
    .CK(clknet_3_4__leaf_clk),
    .Q(prodm3_s1[0]),
    .QN(_043_));
 DFF_X1 _153_ (.D(prodm3_s0[1]),
    .CK(clknet_3_3__leaf_clk),
    .Q(prodm3_s1[1]),
    .QN(_042_));
 DFF_X1 _154_ (.D(prodm3_s0[2]),
    .CK(clknet_3_3__leaf_clk),
    .Q(prodm3_s1[2]),
    .QN(_041_));
 DFF_X1 _155_ (.D(prodm3_s0[3]),
    .CK(clknet_3_1__leaf_clk),
    .Q(prodm3_s1[3]),
    .QN(_040_));
 DFF_X1 _156_ (.D(prodm3_s0[4]),
    .CK(clknet_3_0__leaf_clk),
    .Q(prodm3_s1[4]),
    .QN(_039_));
 DFF_X1 _157_ (.D(prodm3_s0[5]),
    .CK(clknet_3_0__leaf_clk),
    .Q(prodm3_s1[5]),
    .QN(_038_));
 DFF_X1 _158_ (.D(prodm3_s0[6]),
    .CK(clknet_3_0__leaf_clk),
    .Q(prodm3_s1[6]),
    .QN(_037_));
 DFF_X1 _159_ (.D(prodm3_s0[7]),
    .CK(clknet_3_0__leaf_clk),
    .Q(prodm3_s1[7]),
    .QN(_095_));
 DFF_X1 _160_ (.D(sums1[0]),
    .CK(clknet_3_5__leaf_clk),
    .Q(sum_s1[0]),
    .QN(_036_));
 DFF_X2 _161_ (.D(sums1[1]),
    .CK(clknet_3_4__leaf_clk),
    .Q(sum_s1[1]),
    .QN(_035_));
 DFF_X2 _162_ (.D(sums1[2]),
    .CK(clknet_3_7__leaf_clk),
    .Q(sum_s1[2]),
    .QN(_034_));
 DFF_X2 _163_ (.D(sums1[3]),
    .CK(clknet_3_4__leaf_clk),
    .Q(sum_s1[3]),
    .QN(_033_));
 DFF_X2 _164_ (.D(sums1[4]),
    .CK(clknet_3_3__leaf_clk),
    .Q(sum_s1[4]),
    .QN(_032_));
 DFF_X2 _165_ (.D(sums1[5]),
    .CK(clknet_3_6__leaf_clk),
    .Q(sum_s1[5]),
    .QN(_031_));
 DFF_X2 _166_ (.D(sums1[6]),
    .CK(clknet_3_3__leaf_clk),
    .Q(sum_s1[6]),
    .QN(_030_));
 DFF_X2 _167_ (.D(sums1[7]),
    .CK(clknet_3_3__leaf_clk),
    .Q(sum_s1[7]),
    .QN(_096_));
 DFF_X1 _168_ (.D(prodm0[0]),
    .CK(clknet_3_6__leaf_clk),
    .Q(prodm0_s0[0]),
    .QN(_029_));
 DFF_X1 _169_ (.D(prodm0[1]),
    .CK(clknet_3_0__leaf_clk),
    .Q(prodm0_s0[1]),
    .QN(_028_));
 DFF_X1 _170_ (.D(prodm0[2]),
    .CK(clknet_3_7__leaf_clk),
    .Q(prodm0_s0[2]),
    .QN(_027_));
 DFF_X1 _171_ (.D(prodm0[3]),
    .CK(clknet_3_7__leaf_clk),
    .Q(prodm0_s0[3]),
    .QN(_026_));
 DFF_X1 _172_ (.D(prodm0[4]),
    .CK(clknet_3_5__leaf_clk),
    .Q(prodm0_s0[4]),
    .QN(_025_));
 DFF_X1 _173_ (.D(prodm0[5]),
    .CK(clknet_3_5__leaf_clk),
    .Q(prodm0_s0[5]),
    .QN(_024_));
 DFF_X1 _174_ (.D(prodm0[6]),
    .CK(clknet_3_5__leaf_clk),
    .Q(prodm0_s0[6]),
    .QN(_023_));
 DFF_X1 _175_ (.D(prodm0[7]),
    .CK(clknet_3_6__leaf_clk),
    .Q(prodm0_s0[7]),
    .QN(_097_));
 DFF_X2 _176_ (.D(prodm1[0]),
    .CK(clknet_3_4__leaf_clk),
    .Q(prodm1_s0[0]),
    .QN(_022_));
 DFF_X2 _177_ (.D(prodm1[1]),
    .CK(clknet_3_5__leaf_clk),
    .Q(prodm1_s0[1]),
    .QN(_021_));
 DFF_X2 _178_ (.D(prodm1[2]),
    .CK(clknet_3_4__leaf_clk),
    .Q(prodm1_s0[2]),
    .QN(_020_));
 DFF_X2 _179_ (.D(prodm1[3]),
    .CK(clknet_3_4__leaf_clk),
    .Q(prodm1_s0[3]),
    .QN(_019_));
 DFF_X2 _180_ (.D(prodm1[4]),
    .CK(clknet_3_1__leaf_clk),
    .Q(prodm1_s0[4]),
    .QN(_018_));
 DFF_X2 _181_ (.D(prodm1[5]),
    .CK(clknet_3_1__leaf_clk),
    .Q(prodm1_s0[5]),
    .QN(_017_));
 DFF_X2 _182_ (.D(prodm1[6]),
    .CK(clknet_3_1__leaf_clk),
    .Q(prodm1_s0[6]),
    .QN(_016_));
 DFF_X2 _183_ (.D(prodm1[7]),
    .CK(clknet_3_1__leaf_clk),
    .Q(prodm1_s0[7]),
    .QN(_098_));
 DFF_X2 _184_ (.D(prodm2[0]),
    .CK(clknet_3_4__leaf_clk),
    .Q(prodm2_s0[0]),
    .QN(_015_));
 DFF_X2 _185_ (.D(prodm2[1]),
    .CK(clknet_3_1__leaf_clk),
    .Q(prodm2_s0[1]),
    .QN(_014_));
 DFF_X2 _186_ (.D(prodm2[2]),
    .CK(clknet_3_2__leaf_clk),
    .Q(prodm2_s0[2]),
    .QN(_013_));
 DFF_X2 _187_ (.D(prodm2[3]),
    .CK(clknet_3_1__leaf_clk),
    .Q(prodm2_s0[3]),
    .QN(_012_));
 DFF_X2 _188_ (.D(prodm2[4]),
    .CK(clknet_3_2__leaf_clk),
    .Q(prodm2_s0[4]),
    .QN(_011_));
 DFF_X2 _189_ (.D(prodm2[5]),
    .CK(clknet_3_3__leaf_clk),
    .Q(prodm2_s0[5]),
    .QN(_010_));
 DFF_X2 _190_ (.D(prodm2[6]),
    .CK(clknet_3_2__leaf_clk),
    .Q(prodm2_s0[6]),
    .QN(_009_));
 DFF_X2 _191_ (.D(prodm2[7]),
    .CK(clknet_3_3__leaf_clk),
    .Q(prodm2_s0[7]),
    .QN(_099_));
 DFF_X1 _192_ (.D(prodm3[0]),
    .CK(clknet_3_4__leaf_clk),
    .Q(prodm3_s0[0]),
    .QN(_008_));
 DFF_X1 _193_ (.D(prodm3[1]),
    .CK(clknet_3_1__leaf_clk),
    .Q(prodm3_s0[1]),
    .QN(_007_));
 DFF_X1 _194_ (.D(prodm3[2]),
    .CK(clknet_3_1__leaf_clk),
    .Q(prodm3_s0[2]),
    .QN(_006_));
 DFF_X1 _195_ (.D(prodm3[3]),
    .CK(clknet_3_1__leaf_clk),
    .Q(prodm3_s0[3]),
    .QN(_005_));
 DFF_X1 _196_ (.D(prodm3[4]),
    .CK(clknet_3_0__leaf_clk),
    .Q(prodm3_s0[4]),
    .QN(_004_));
 DFF_X1 _197_ (.D(prodm3[5]),
    .CK(clknet_3_0__leaf_clk),
    .Q(prodm3_s0[5]),
    .QN(_003_));
 DFF_X1 _198_ (.D(prodm3[6]),
    .CK(clknet_3_0__leaf_clk),
    .Q(prodm3_s0[6]),
    .QN(_002_));
 DFF_X1 _199_ (.D(prodm3[7]),
    .CK(clknet_3_0__leaf_clk),
    .Q(prodm3_s0[7]),
    .QN(_001_));
 AND2_X1 \stage1/FA1_0/HA1/_0_  (.A1(prodm1_s0[0]),
    .A2(prodm2_s0[0]),
    .ZN(\stage1/FA1_0/ha1_carry ));
 XOR2_X2 \stage1/FA1_0/HA1/_1_  (.A(prodm1_s0[0]),
    .B(prodm2_s0[0]),
    .Z(\stage1/FA1_0/ha1_sum ));
 AND2_X1 \stage1/FA1_0/HA2/_0_  (.A1(\stage1/FA1_0/ha1_sum ),
    .A2(\stage1/_07_ ),
    .ZN(\stage1/FA1_0/ha2_carry ));
 XOR2_X1 \stage1/FA1_0/HA2/_1_  (.A(\stage1/FA1_0/ha1_sum ),
    .B(\stage1/_07_ ),
    .Z(\stage1/sum1 [0]));
 OR2_X1 \stage1/FA1_0/_0_  (.A1(\stage1/FA1_0/ha1_carry ),
    .A2(\stage1/FA1_0/ha2_carry ),
    .ZN(\stage1/carry1 [0]));
 AND2_X1 \stage1/HA0_0/_0_  (.A1(prodm1_s0[0]),
    .A2(prodm2_s0[0]),
    .ZN(\stage1/carry0 [0]));
 XOR2_X1 \stage1/HA0_0/_1_  (.A(prodm1_s0[0]),
    .B(prodm2_s0[0]),
    .Z(\stage1/sum0 [0]));
 INV_X4 \stage1/_08_  (.A(ground),
    .ZN(\stage1/_07_ ));
 MUX2_X1 \stage1/_09_  (.A(\stage1/sum0 [0]),
    .B(\stage1/sum1 [0]),
    .S(ground),
    .Z(sums1[0]));
 MUX2_X1 \stage1/_10_  (.A(\stage1/carry0 [0]),
    .B(\stage1/carry1 [0]),
    .S(ground),
    .Z(\stage1/_00_ ));
 MUX2_X1 \stage1/_11_  (.A(\stage1/sum0 [1]),
    .B(\stage1/sum1 [1]),
    .S(\stage1/_00_ ),
    .Z(sums1[1]));
 MUX2_X1 \stage1/_12_  (.A(\stage1/carry0 [1]),
    .B(\stage1/carry1 [1]),
    .S(\stage1/_00_ ),
    .Z(\stage1/_01_ ));
 MUX2_X1 \stage1/_13_  (.A(\stage1/sum0 [2]),
    .B(\stage1/sum1 [2]),
    .S(\stage1/_01_ ),
    .Z(sums1[2]));
 MUX2_X1 \stage1/_14_  (.A(\stage1/carry0 [2]),
    .B(\stage1/carry1 [2]),
    .S(\stage1/_01_ ),
    .Z(\stage1/_02_ ));
 MUX2_X1 \stage1/_15_  (.A(\stage1/sum0 [3]),
    .B(\stage1/sum1 [3]),
    .S(\stage1/_02_ ),
    .Z(sums1[3]));
 MUX2_X1 \stage1/_16_  (.A(\stage1/carry0 [3]),
    .B(\stage1/carry1 [3]),
    .S(\stage1/_02_ ),
    .Z(\stage1/_03_ ));
 MUX2_X1 \stage1/_17_  (.A(\stage1/sum0 [4]),
    .B(\stage1/sum1 [4]),
    .S(\stage1/_03_ ),
    .Z(sums1[4]));
 MUX2_X1 \stage1/_18_  (.A(\stage1/carry0 [4]),
    .B(\stage1/carry1 [4]),
    .S(\stage1/_03_ ),
    .Z(\stage1/_04_ ));
 MUX2_X1 \stage1/_19_  (.A(\stage1/sum0 [5]),
    .B(\stage1/sum1 [5]),
    .S(\stage1/_04_ ),
    .Z(sums1[5]));
 MUX2_X1 \stage1/_20_  (.A(\stage1/carry0 [5]),
    .B(\stage1/carry1 [5]),
    .S(\stage1/_04_ ),
    .Z(\stage1/_05_ ));
 MUX2_X1 \stage1/_21_  (.A(\stage1/sum0 [6]),
    .B(\stage1/sum1 [6]),
    .S(\stage1/_05_ ),
    .Z(sums1[6]));
 MUX2_X1 \stage1/_22_  (.A(\stage1/carry0 [6]),
    .B(\stage1/carry1 [6]),
    .S(\stage1/_05_ ),
    .Z(\stage1/_06_ ));
 MUX2_X1 \stage1/_23_  (.A(\stage1/sum0 [7]),
    .B(\stage1/sum1 [7]),
    .S(\stage1/_06_ ),
    .Z(sums1[7]));
 MUX2_X1 \stage1/_24_  (.A(\stage1/carry0 [7]),
    .B(\stage1/carry1 [7]),
    .S(\stage1/_06_ ),
    .Z(c1));
 AND2_X1 \stage1/gen_csa[1].FA0/HA1/_0_  (.A1(prodm1_s0[1]),
    .A2(prodm2_s0[1]),
    .ZN(\stage1/gen_csa[1].FA0/ha1_carry ));
 XOR2_X2 \stage1/gen_csa[1].FA0/HA1/_1_  (.A(prodm1_s0[1]),
    .B(prodm2_s0[1]),
    .Z(\stage1/gen_csa[1].FA0/ha1_sum ));
 AND2_X1 \stage1/gen_csa[1].FA0/HA2/_0_  (.A1(\stage1/gen_csa[1].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\stage1/gen_csa[1].FA0/ha2_carry ));
 XOR2_X1 \stage1/gen_csa[1].FA0/HA2/_1_  (.A(\stage1/gen_csa[1].FA0/ha1_sum ),
    .B(ground),
    .Z(\stage1/sum0 [1]));
 OR2_X1 \stage1/gen_csa[1].FA0/_0_  (.A1(\stage1/gen_csa[1].FA0/ha1_carry ),
    .A2(\stage1/gen_csa[1].FA0/ha2_carry ),
    .ZN(\stage1/carry0 [1]));
 AND2_X1 \stage1/gen_csa[1].FA1/HA1/_0_  (.A1(prodm1_s0[1]),
    .A2(prodm2_s0[1]),
    .ZN(\stage1/gen_csa[1].FA1/ha1_carry ));
 XOR2_X2 \stage1/gen_csa[1].FA1/HA1/_1_  (.A(prodm1_s0[1]),
    .B(prodm2_s0[1]),
    .Z(\stage1/gen_csa[1].FA1/ha1_sum ));
 AND2_X1 \stage1/gen_csa[1].FA1/HA2/_0_  (.A1(\stage1/gen_csa[1].FA1/ha1_sum ),
    .A2(\stage1/_07_ ),
    .ZN(\stage1/gen_csa[1].FA1/ha2_carry ));
 XOR2_X1 \stage1/gen_csa[1].FA1/HA2/_1_  (.A(\stage1/gen_csa[1].FA1/ha1_sum ),
    .B(\stage1/_07_ ),
    .Z(\stage1/sum1 [1]));
 OR2_X1 \stage1/gen_csa[1].FA1/_0_  (.A1(\stage1/gen_csa[1].FA1/ha1_carry ),
    .A2(\stage1/gen_csa[1].FA1/ha2_carry ),
    .ZN(\stage1/carry1 [1]));
 AND2_X1 \stage1/gen_csa[2].FA0/HA1/_0_  (.A1(prodm1_s0[2]),
    .A2(prodm2_s0[2]),
    .ZN(\stage1/gen_csa[2].FA0/ha1_carry ));
 XOR2_X2 \stage1/gen_csa[2].FA0/HA1/_1_  (.A(prodm1_s0[2]),
    .B(prodm2_s0[2]),
    .Z(\stage1/gen_csa[2].FA0/ha1_sum ));
 AND2_X1 \stage1/gen_csa[2].FA0/HA2/_0_  (.A1(\stage1/gen_csa[2].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\stage1/gen_csa[2].FA0/ha2_carry ));
 XOR2_X1 \stage1/gen_csa[2].FA0/HA2/_1_  (.A(\stage1/gen_csa[2].FA0/ha1_sum ),
    .B(ground),
    .Z(\stage1/sum0 [2]));
 OR2_X1 \stage1/gen_csa[2].FA0/_0_  (.A1(\stage1/gen_csa[2].FA0/ha1_carry ),
    .A2(\stage1/gen_csa[2].FA0/ha2_carry ),
    .ZN(\stage1/carry0 [2]));
 AND2_X1 \stage1/gen_csa[2].FA1/HA1/_0_  (.A1(prodm1_s0[2]),
    .A2(prodm2_s0[2]),
    .ZN(\stage1/gen_csa[2].FA1/ha1_carry ));
 XOR2_X2 \stage1/gen_csa[2].FA1/HA1/_1_  (.A(prodm1_s0[2]),
    .B(prodm2_s0[2]),
    .Z(\stage1/gen_csa[2].FA1/ha1_sum ));
 AND2_X1 \stage1/gen_csa[2].FA1/HA2/_0_  (.A1(\stage1/gen_csa[2].FA1/ha1_sum ),
    .A2(\stage1/_07_ ),
    .ZN(\stage1/gen_csa[2].FA1/ha2_carry ));
 XOR2_X1 \stage1/gen_csa[2].FA1/HA2/_1_  (.A(\stage1/gen_csa[2].FA1/ha1_sum ),
    .B(\stage1/_07_ ),
    .Z(\stage1/sum1 [2]));
 OR2_X1 \stage1/gen_csa[2].FA1/_0_  (.A1(\stage1/gen_csa[2].FA1/ha1_carry ),
    .A2(\stage1/gen_csa[2].FA1/ha2_carry ),
    .ZN(\stage1/carry1 [2]));
 AND2_X1 \stage1/gen_csa[3].FA0/HA1/_0_  (.A1(prodm1_s0[3]),
    .A2(prodm2_s0[3]),
    .ZN(\stage1/gen_csa[3].FA0/ha1_carry ));
 XOR2_X2 \stage1/gen_csa[3].FA0/HA1/_1_  (.A(prodm1_s0[3]),
    .B(prodm2_s0[3]),
    .Z(\stage1/gen_csa[3].FA0/ha1_sum ));
 AND2_X1 \stage1/gen_csa[3].FA0/HA2/_0_  (.A1(\stage1/gen_csa[3].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\stage1/gen_csa[3].FA0/ha2_carry ));
 XOR2_X1 \stage1/gen_csa[3].FA0/HA2/_1_  (.A(\stage1/gen_csa[3].FA0/ha1_sum ),
    .B(ground),
    .Z(\stage1/sum0 [3]));
 OR2_X1 \stage1/gen_csa[3].FA0/_0_  (.A1(\stage1/gen_csa[3].FA0/ha1_carry ),
    .A2(\stage1/gen_csa[3].FA0/ha2_carry ),
    .ZN(\stage1/carry0 [3]));
 AND2_X1 \stage1/gen_csa[3].FA1/HA1/_0_  (.A1(prodm1_s0[3]),
    .A2(prodm2_s0[3]),
    .ZN(\stage1/gen_csa[3].FA1/ha1_carry ));
 XOR2_X2 \stage1/gen_csa[3].FA1/HA1/_1_  (.A(prodm1_s0[3]),
    .B(prodm2_s0[3]),
    .Z(\stage1/gen_csa[3].FA1/ha1_sum ));
 AND2_X1 \stage1/gen_csa[3].FA1/HA2/_0_  (.A1(\stage1/gen_csa[3].FA1/ha1_sum ),
    .A2(\stage1/_07_ ),
    .ZN(\stage1/gen_csa[3].FA1/ha2_carry ));
 XOR2_X1 \stage1/gen_csa[3].FA1/HA2/_1_  (.A(\stage1/gen_csa[3].FA1/ha1_sum ),
    .B(\stage1/_07_ ),
    .Z(\stage1/sum1 [3]));
 OR2_X1 \stage1/gen_csa[3].FA1/_0_  (.A1(\stage1/gen_csa[3].FA1/ha1_carry ),
    .A2(\stage1/gen_csa[3].FA1/ha2_carry ),
    .ZN(\stage1/carry1 [3]));
 AND2_X1 \stage1/gen_csa[4].FA0/HA1/_0_  (.A1(prodm1_s0[4]),
    .A2(prodm2_s0[4]),
    .ZN(\stage1/gen_csa[4].FA0/ha1_carry ));
 XOR2_X2 \stage1/gen_csa[4].FA0/HA1/_1_  (.A(prodm1_s0[4]),
    .B(prodm2_s0[4]),
    .Z(\stage1/gen_csa[4].FA0/ha1_sum ));
 AND2_X1 \stage1/gen_csa[4].FA0/HA2/_0_  (.A1(\stage1/gen_csa[4].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\stage1/gen_csa[4].FA0/ha2_carry ));
 XOR2_X1 \stage1/gen_csa[4].FA0/HA2/_1_  (.A(\stage1/gen_csa[4].FA0/ha1_sum ),
    .B(ground),
    .Z(\stage1/sum0 [4]));
 OR2_X1 \stage1/gen_csa[4].FA0/_0_  (.A1(\stage1/gen_csa[4].FA0/ha1_carry ),
    .A2(\stage1/gen_csa[4].FA0/ha2_carry ),
    .ZN(\stage1/carry0 [4]));
 AND2_X1 \stage1/gen_csa[4].FA1/HA1/_0_  (.A1(prodm1_s0[4]),
    .A2(prodm2_s0[4]),
    .ZN(\stage1/gen_csa[4].FA1/ha1_carry ));
 XOR2_X2 \stage1/gen_csa[4].FA1/HA1/_1_  (.A(prodm1_s0[4]),
    .B(prodm2_s0[4]),
    .Z(\stage1/gen_csa[4].FA1/ha1_sum ));
 AND2_X1 \stage1/gen_csa[4].FA1/HA2/_0_  (.A1(\stage1/gen_csa[4].FA1/ha1_sum ),
    .A2(\stage1/_07_ ),
    .ZN(\stage1/gen_csa[4].FA1/ha2_carry ));
 XOR2_X1 \stage1/gen_csa[4].FA1/HA2/_1_  (.A(\stage1/gen_csa[4].FA1/ha1_sum ),
    .B(\stage1/_07_ ),
    .Z(\stage1/sum1 [4]));
 OR2_X1 \stage1/gen_csa[4].FA1/_0_  (.A1(\stage1/gen_csa[4].FA1/ha1_carry ),
    .A2(\stage1/gen_csa[4].FA1/ha2_carry ),
    .ZN(\stage1/carry1 [4]));
 AND2_X1 \stage1/gen_csa[5].FA0/HA1/_0_  (.A1(prodm1_s0[5]),
    .A2(prodm2_s0[5]),
    .ZN(\stage1/gen_csa[5].FA0/ha1_carry ));
 XOR2_X2 \stage1/gen_csa[5].FA0/HA1/_1_  (.A(prodm1_s0[5]),
    .B(prodm2_s0[5]),
    .Z(\stage1/gen_csa[5].FA0/ha1_sum ));
 AND2_X1 \stage1/gen_csa[5].FA0/HA2/_0_  (.A1(\stage1/gen_csa[5].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\stage1/gen_csa[5].FA0/ha2_carry ));
 XOR2_X1 \stage1/gen_csa[5].FA0/HA2/_1_  (.A(\stage1/gen_csa[5].FA0/ha1_sum ),
    .B(ground),
    .Z(\stage1/sum0 [5]));
 OR2_X1 \stage1/gen_csa[5].FA0/_0_  (.A1(\stage1/gen_csa[5].FA0/ha1_carry ),
    .A2(\stage1/gen_csa[5].FA0/ha2_carry ),
    .ZN(\stage1/carry0 [5]));
 AND2_X1 \stage1/gen_csa[5].FA1/HA1/_0_  (.A1(prodm1_s0[5]),
    .A2(prodm2_s0[5]),
    .ZN(\stage1/gen_csa[5].FA1/ha1_carry ));
 XOR2_X1 \stage1/gen_csa[5].FA1/HA1/_1_  (.A(prodm1_s0[5]),
    .B(prodm2_s0[5]),
    .Z(\stage1/gen_csa[5].FA1/ha1_sum ));
 AND2_X1 \stage1/gen_csa[5].FA1/HA2/_0_  (.A1(\stage1/gen_csa[5].FA1/ha1_sum ),
    .A2(\stage1/_07_ ),
    .ZN(\stage1/gen_csa[5].FA1/ha2_carry ));
 XOR2_X1 \stage1/gen_csa[5].FA1/HA2/_1_  (.A(\stage1/gen_csa[5].FA1/ha1_sum ),
    .B(\stage1/_07_ ),
    .Z(\stage1/sum1 [5]));
 OR2_X1 \stage1/gen_csa[5].FA1/_0_  (.A1(\stage1/gen_csa[5].FA1/ha1_carry ),
    .A2(\stage1/gen_csa[5].FA1/ha2_carry ),
    .ZN(\stage1/carry1 [5]));
 AND2_X1 \stage1/gen_csa[6].FA0/HA1/_0_  (.A1(prodm1_s0[6]),
    .A2(prodm2_s0[6]),
    .ZN(\stage1/gen_csa[6].FA0/ha1_carry ));
 XOR2_X2 \stage1/gen_csa[6].FA0/HA1/_1_  (.A(prodm1_s0[6]),
    .B(prodm2_s0[6]),
    .Z(\stage1/gen_csa[6].FA0/ha1_sum ));
 AND2_X1 \stage1/gen_csa[6].FA0/HA2/_0_  (.A1(\stage1/gen_csa[6].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\stage1/gen_csa[6].FA0/ha2_carry ));
 XOR2_X1 \stage1/gen_csa[6].FA0/HA2/_1_  (.A(\stage1/gen_csa[6].FA0/ha1_sum ),
    .B(ground),
    .Z(\stage1/sum0 [6]));
 OR2_X1 \stage1/gen_csa[6].FA0/_0_  (.A1(\stage1/gen_csa[6].FA0/ha1_carry ),
    .A2(\stage1/gen_csa[6].FA0/ha2_carry ),
    .ZN(\stage1/carry0 [6]));
 AND2_X1 \stage1/gen_csa[6].FA1/HA1/_0_  (.A1(prodm1_s0[6]),
    .A2(prodm2_s0[6]),
    .ZN(\stage1/gen_csa[6].FA1/ha1_carry ));
 XOR2_X2 \stage1/gen_csa[6].FA1/HA1/_1_  (.A(prodm1_s0[6]),
    .B(prodm2_s0[6]),
    .Z(\stage1/gen_csa[6].FA1/ha1_sum ));
 AND2_X1 \stage1/gen_csa[6].FA1/HA2/_0_  (.A1(\stage1/gen_csa[6].FA1/ha1_sum ),
    .A2(\stage1/_07_ ),
    .ZN(\stage1/gen_csa[6].FA1/ha2_carry ));
 XOR2_X1 \stage1/gen_csa[6].FA1/HA2/_1_  (.A(\stage1/gen_csa[6].FA1/ha1_sum ),
    .B(\stage1/_07_ ),
    .Z(\stage1/sum1 [6]));
 OR2_X1 \stage1/gen_csa[6].FA1/_0_  (.A1(\stage1/gen_csa[6].FA1/ha1_carry ),
    .A2(\stage1/gen_csa[6].FA1/ha2_carry ),
    .ZN(\stage1/carry1 [6]));
 AND2_X1 \stage1/gen_csa[7].FA0/HA1/_0_  (.A1(prodm1_s0[7]),
    .A2(prodm2_s0[7]),
    .ZN(\stage1/gen_csa[7].FA0/ha1_carry ));
 XOR2_X2 \stage1/gen_csa[7].FA0/HA1/_1_  (.A(prodm1_s0[7]),
    .B(prodm2_s0[7]),
    .Z(\stage1/gen_csa[7].FA0/ha1_sum ));
 AND2_X1 \stage1/gen_csa[7].FA0/HA2/_0_  (.A1(\stage1/gen_csa[7].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\stage1/gen_csa[7].FA0/ha2_carry ));
 XOR2_X1 \stage1/gen_csa[7].FA0/HA2/_1_  (.A(\stage1/gen_csa[7].FA0/ha1_sum ),
    .B(ground),
    .Z(\stage1/sum0 [7]));
 OR2_X1 \stage1/gen_csa[7].FA0/_0_  (.A1(\stage1/gen_csa[7].FA0/ha1_carry ),
    .A2(\stage1/gen_csa[7].FA0/ha2_carry ),
    .ZN(\stage1/carry0 [7]));
 AND2_X1 \stage1/gen_csa[7].FA1/HA1/_0_  (.A1(prodm1_s0[7]),
    .A2(prodm2_s0[7]),
    .ZN(\stage1/gen_csa[7].FA1/ha1_carry ));
 XOR2_X2 \stage1/gen_csa[7].FA1/HA1/_1_  (.A(prodm1_s0[7]),
    .B(prodm2_s0[7]),
    .Z(\stage1/gen_csa[7].FA1/ha1_sum ));
 AND2_X1 \stage1/gen_csa[7].FA1/HA2/_0_  (.A1(\stage1/gen_csa[7].FA1/ha1_sum ),
    .A2(\stage1/_07_ ),
    .ZN(\stage1/gen_csa[7].FA1/ha2_carry ));
 XOR2_X1 \stage1/gen_csa[7].FA1/HA2/_1_  (.A(\stage1/gen_csa[7].FA1/ha1_sum ),
    .B(\stage1/_07_ ),
    .Z(\stage1/sum1 [7]));
 OR2_X1 \stage1/gen_csa[7].FA1/_0_  (.A1(\stage1/gen_csa[7].FA1/ha1_carry ),
    .A2(\stage1/gen_csa[7].FA1/ha2_carry ),
    .ZN(\stage1/carry1 [7]));
 AND2_X1 \stage2/FA1_0/HA1/_0_  (.A1(prodm0_s1[4]),
    .A2(sum_s1[0]),
    .ZN(\stage2/FA1_0/ha1_carry ));
 XOR2_X1 \stage2/FA1_0/HA1/_1_  (.A(prodm0_s1[4]),
    .B(sum_s1[0]),
    .Z(\stage2/FA1_0/ha1_sum ));
 AND2_X1 \stage2/FA1_0/HA2/_0_  (.A1(\stage2/FA1_0/ha1_sum ),
    .A2(\stage2/_07_ ),
    .ZN(\stage2/FA1_0/ha2_carry ));
 XOR2_X1 \stage2/FA1_0/HA2/_1_  (.A(\stage2/FA1_0/ha1_sum ),
    .B(\stage2/_07_ ),
    .Z(\stage2/sum1 [0]));
 OR2_X1 \stage2/FA1_0/_0_  (.A1(\stage2/FA1_0/ha1_carry ),
    .A2(\stage2/FA1_0/ha2_carry ),
    .ZN(\stage2/carry1 [0]));
 AND2_X1 \stage2/HA0_0/_0_  (.A1(prodm0_s1[4]),
    .A2(sum_s1[0]),
    .ZN(\stage2/carry0 [0]));
 XOR2_X1 \stage2/HA0_0/_1_  (.A(prodm0_s1[4]),
    .B(sum_s1[0]),
    .Z(\stage2/sum0 [0]));
 INV_X4 \stage2/_08_  (.A(ground),
    .ZN(\stage2/_07_ ));
 MUX2_X1 \stage2/_09_  (.A(\stage2/sum0 [0]),
    .B(\stage2/sum1 [0]),
    .S(ground),
    .Z(sums2[0]));
 MUX2_X1 \stage2/_10_  (.A(\stage2/carry0 [0]),
    .B(\stage2/carry1 [0]),
    .S(ground),
    .Z(\stage2/_00_ ));
 MUX2_X1 \stage2/_11_  (.A(\stage2/sum0 [1]),
    .B(\stage2/sum1 [1]),
    .S(\stage2/_00_ ),
    .Z(sums2[1]));
 MUX2_X1 \stage2/_12_  (.A(\stage2/carry0 [1]),
    .B(\stage2/carry1 [1]),
    .S(\stage2/_00_ ),
    .Z(\stage2/_01_ ));
 MUX2_X1 \stage2/_13_  (.A(\stage2/sum0 [2]),
    .B(\stage2/sum1 [2]),
    .S(\stage2/_01_ ),
    .Z(sums2[2]));
 MUX2_X1 \stage2/_14_  (.A(\stage2/carry0 [2]),
    .B(\stage2/carry1 [2]),
    .S(\stage2/_01_ ),
    .Z(\stage2/_02_ ));
 MUX2_X1 \stage2/_15_  (.A(\stage2/sum0 [3]),
    .B(\stage2/sum1 [3]),
    .S(\stage2/_02_ ),
    .Z(sums2[3]));
 MUX2_X1 \stage2/_16_  (.A(\stage2/carry0 [3]),
    .B(\stage2/carry1 [3]),
    .S(\stage2/_02_ ),
    .Z(\stage2/_03_ ));
 MUX2_X1 \stage2/_17_  (.A(\stage2/sum0 [4]),
    .B(\stage2/sum1 [4]),
    .S(\stage2/_03_ ),
    .Z(sums2[4]));
 MUX2_X1 \stage2/_18_  (.A(\stage2/carry0 [4]),
    .B(\stage2/carry1 [4]),
    .S(\stage2/_03_ ),
    .Z(\stage2/_04_ ));
 MUX2_X1 \stage2/_19_  (.A(\stage2/sum0 [5]),
    .B(\stage2/sum1 [5]),
    .S(\stage2/_04_ ),
    .Z(sums2[5]));
 MUX2_X1 \stage2/_20_  (.A(\stage2/carry0 [5]),
    .B(\stage2/carry1 [5]),
    .S(\stage2/_04_ ),
    .Z(\stage2/_05_ ));
 MUX2_X1 \stage2/_21_  (.A(\stage2/sum0 [6]),
    .B(\stage2/sum1 [6]),
    .S(\stage2/_05_ ),
    .Z(sums2[6]));
 MUX2_X1 \stage2/_22_  (.A(\stage2/carry0 [6]),
    .B(\stage2/carry1 [6]),
    .S(\stage2/_05_ ),
    .Z(\stage2/_06_ ));
 MUX2_X1 \stage2/_23_  (.A(\stage2/sum0 [7]),
    .B(\stage2/sum1 [7]),
    .S(\stage2/_06_ ),
    .Z(sums2[7]));
 MUX2_X1 \stage2/_24_  (.A(\stage2/carry0 [7]),
    .B(\stage2/carry1 [7]),
    .S(\stage2/_06_ ),
    .Z(c2));
 AND2_X1 \stage2/gen_csa[1].FA0/HA1/_0_  (.A1(prodm0_s1[5]),
    .A2(sum_s1[1]),
    .ZN(\stage2/gen_csa[1].FA0/ha1_carry ));
 XOR2_X2 \stage2/gen_csa[1].FA0/HA1/_1_  (.A(prodm0_s1[5]),
    .B(sum_s1[1]),
    .Z(\stage2/gen_csa[1].FA0/ha1_sum ));
 AND2_X1 \stage2/gen_csa[1].FA0/HA2/_0_  (.A1(\stage2/gen_csa[1].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\stage2/gen_csa[1].FA0/ha2_carry ));
 XOR2_X1 \stage2/gen_csa[1].FA0/HA2/_1_  (.A(\stage2/gen_csa[1].FA0/ha1_sum ),
    .B(ground),
    .Z(\stage2/sum0 [1]));
 OR2_X1 \stage2/gen_csa[1].FA0/_0_  (.A1(\stage2/gen_csa[1].FA0/ha1_carry ),
    .A2(\stage2/gen_csa[1].FA0/ha2_carry ),
    .ZN(\stage2/carry0 [1]));
 AND2_X1 \stage2/gen_csa[1].FA1/HA1/_0_  (.A1(prodm0_s1[5]),
    .A2(sum_s1[1]),
    .ZN(\stage2/gen_csa[1].FA1/ha1_carry ));
 XOR2_X2 \stage2/gen_csa[1].FA1/HA1/_1_  (.A(prodm0_s1[5]),
    .B(sum_s1[1]),
    .Z(\stage2/gen_csa[1].FA1/ha1_sum ));
 AND2_X1 \stage2/gen_csa[1].FA1/HA2/_0_  (.A1(\stage2/gen_csa[1].FA1/ha1_sum ),
    .A2(\stage2/_07_ ),
    .ZN(\stage2/gen_csa[1].FA1/ha2_carry ));
 XOR2_X1 \stage2/gen_csa[1].FA1/HA2/_1_  (.A(\stage2/gen_csa[1].FA1/ha1_sum ),
    .B(\stage2/_07_ ),
    .Z(\stage2/sum1 [1]));
 OR2_X1 \stage2/gen_csa[1].FA1/_0_  (.A1(\stage2/gen_csa[1].FA1/ha1_carry ),
    .A2(\stage2/gen_csa[1].FA1/ha2_carry ),
    .ZN(\stage2/carry1 [1]));
 AND2_X1 \stage2/gen_csa[2].FA0/HA1/_0_  (.A1(prodm0_s1[6]),
    .A2(sum_s1[2]),
    .ZN(\stage2/gen_csa[2].FA0/ha1_carry ));
 XOR2_X2 \stage2/gen_csa[2].FA0/HA1/_1_  (.A(prodm0_s1[6]),
    .B(sum_s1[2]),
    .Z(\stage2/gen_csa[2].FA0/ha1_sum ));
 AND2_X1 \stage2/gen_csa[2].FA0/HA2/_0_  (.A1(\stage2/gen_csa[2].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\stage2/gen_csa[2].FA0/ha2_carry ));
 XOR2_X1 \stage2/gen_csa[2].FA0/HA2/_1_  (.A(\stage2/gen_csa[2].FA0/ha1_sum ),
    .B(ground),
    .Z(\stage2/sum0 [2]));
 OR2_X1 \stage2/gen_csa[2].FA0/_0_  (.A1(\stage2/gen_csa[2].FA0/ha1_carry ),
    .A2(\stage2/gen_csa[2].FA0/ha2_carry ),
    .ZN(\stage2/carry0 [2]));
 AND2_X1 \stage2/gen_csa[2].FA1/HA1/_0_  (.A1(prodm0_s1[6]),
    .A2(sum_s1[2]),
    .ZN(\stage2/gen_csa[2].FA1/ha1_carry ));
 XOR2_X2 \stage2/gen_csa[2].FA1/HA1/_1_  (.A(prodm0_s1[6]),
    .B(sum_s1[2]),
    .Z(\stage2/gen_csa[2].FA1/ha1_sum ));
 AND2_X1 \stage2/gen_csa[2].FA1/HA2/_0_  (.A1(\stage2/gen_csa[2].FA1/ha1_sum ),
    .A2(\stage2/_07_ ),
    .ZN(\stage2/gen_csa[2].FA1/ha2_carry ));
 XOR2_X1 \stage2/gen_csa[2].FA1/HA2/_1_  (.A(\stage2/gen_csa[2].FA1/ha1_sum ),
    .B(\stage2/_07_ ),
    .Z(\stage2/sum1 [2]));
 OR2_X1 \stage2/gen_csa[2].FA1/_0_  (.A1(\stage2/gen_csa[2].FA1/ha1_carry ),
    .A2(\stage2/gen_csa[2].FA1/ha2_carry ),
    .ZN(\stage2/carry1 [2]));
 AND2_X1 \stage2/gen_csa[3].FA0/HA1/_0_  (.A1(prodm0_s1[7]),
    .A2(sum_s1[3]),
    .ZN(\stage2/gen_csa[3].FA0/ha1_carry ));
 XOR2_X2 \stage2/gen_csa[3].FA0/HA1/_1_  (.A(prodm0_s1[7]),
    .B(sum_s1[3]),
    .Z(\stage2/gen_csa[3].FA0/ha1_sum ));
 AND2_X1 \stage2/gen_csa[3].FA0/HA2/_0_  (.A1(\stage2/gen_csa[3].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\stage2/gen_csa[3].FA0/ha2_carry ));
 XOR2_X1 \stage2/gen_csa[3].FA0/HA2/_1_  (.A(\stage2/gen_csa[3].FA0/ha1_sum ),
    .B(ground),
    .Z(\stage2/sum0 [3]));
 OR2_X1 \stage2/gen_csa[3].FA0/_0_  (.A1(\stage2/gen_csa[3].FA0/ha1_carry ),
    .A2(\stage2/gen_csa[3].FA0/ha2_carry ),
    .ZN(\stage2/carry0 [3]));
 AND2_X1 \stage2/gen_csa[3].FA1/HA1/_0_  (.A1(prodm0_s1[7]),
    .A2(sum_s1[3]),
    .ZN(\stage2/gen_csa[3].FA1/ha1_carry ));
 XOR2_X2 \stage2/gen_csa[3].FA1/HA1/_1_  (.A(prodm0_s1[7]),
    .B(sum_s1[3]),
    .Z(\stage2/gen_csa[3].FA1/ha1_sum ));
 AND2_X1 \stage2/gen_csa[3].FA1/HA2/_0_  (.A1(\stage2/gen_csa[3].FA1/ha1_sum ),
    .A2(\stage2/_07_ ),
    .ZN(\stage2/gen_csa[3].FA1/ha2_carry ));
 XOR2_X1 \stage2/gen_csa[3].FA1/HA2/_1_  (.A(\stage2/gen_csa[3].FA1/ha1_sum ),
    .B(\stage2/_07_ ),
    .Z(\stage2/sum1 [3]));
 OR2_X1 \stage2/gen_csa[3].FA1/_0_  (.A1(\stage2/gen_csa[3].FA1/ha1_carry ),
    .A2(\stage2/gen_csa[3].FA1/ha2_carry ),
    .ZN(\stage2/carry1 [3]));
 AND2_X1 \stage2/gen_csa[4].FA0/HA1/_0_  (.A1(ground),
    .A2(sum_s1[4]),
    .ZN(\stage2/gen_csa[4].FA0/ha1_carry ));
 XOR2_X2 \stage2/gen_csa[4].FA0/HA1/_1_  (.A(ground),
    .B(sum_s1[4]),
    .Z(\stage2/gen_csa[4].FA0/ha1_sum ));
 AND2_X1 \stage2/gen_csa[4].FA0/HA2/_0_  (.A1(\stage2/gen_csa[4].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\stage2/gen_csa[4].FA0/ha2_carry ));
 XOR2_X1 \stage2/gen_csa[4].FA0/HA2/_1_  (.A(\stage2/gen_csa[4].FA0/ha1_sum ),
    .B(ground),
    .Z(\stage2/sum0 [4]));
 OR2_X1 \stage2/gen_csa[4].FA0/_0_  (.A1(\stage2/gen_csa[4].FA0/ha1_carry ),
    .A2(\stage2/gen_csa[4].FA0/ha2_carry ),
    .ZN(\stage2/carry0 [4]));
 AND2_X1 \stage2/gen_csa[4].FA1/HA1/_0_  (.A1(ground),
    .A2(sum_s1[4]),
    .ZN(\stage2/gen_csa[4].FA1/ha1_carry ));
 XOR2_X2 \stage2/gen_csa[4].FA1/HA1/_1_  (.A(ground),
    .B(sum_s1[4]),
    .Z(\stage2/gen_csa[4].FA1/ha1_sum ));
 AND2_X1 \stage2/gen_csa[4].FA1/HA2/_0_  (.A1(\stage2/gen_csa[4].FA1/ha1_sum ),
    .A2(\stage2/_07_ ),
    .ZN(\stage2/gen_csa[4].FA1/ha2_carry ));
 XOR2_X1 \stage2/gen_csa[4].FA1/HA2/_1_  (.A(\stage2/gen_csa[4].FA1/ha1_sum ),
    .B(\stage2/_07_ ),
    .Z(\stage2/sum1 [4]));
 OR2_X1 \stage2/gen_csa[4].FA1/_0_  (.A1(\stage2/gen_csa[4].FA1/ha1_carry ),
    .A2(\stage2/gen_csa[4].FA1/ha2_carry ),
    .ZN(\stage2/carry1 [4]));
 AND2_X1 \stage2/gen_csa[5].FA0/HA1/_0_  (.A1(ground),
    .A2(sum_s1[5]),
    .ZN(\stage2/gen_csa[5].FA0/ha1_carry ));
 XOR2_X2 \stage2/gen_csa[5].FA0/HA1/_1_  (.A(ground),
    .B(sum_s1[5]),
    .Z(\stage2/gen_csa[5].FA0/ha1_sum ));
 AND2_X1 \stage2/gen_csa[5].FA0/HA2/_0_  (.A1(\stage2/gen_csa[5].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\stage2/gen_csa[5].FA0/ha2_carry ));
 XOR2_X1 \stage2/gen_csa[5].FA0/HA2/_1_  (.A(\stage2/gen_csa[5].FA0/ha1_sum ),
    .B(ground),
    .Z(\stage2/sum0 [5]));
 OR2_X1 \stage2/gen_csa[5].FA0/_0_  (.A1(\stage2/gen_csa[5].FA0/ha1_carry ),
    .A2(\stage2/gen_csa[5].FA0/ha2_carry ),
    .ZN(\stage2/carry0 [5]));
 AND2_X1 \stage2/gen_csa[5].FA1/HA1/_0_  (.A1(ground),
    .A2(sum_s1[5]),
    .ZN(\stage2/gen_csa[5].FA1/ha1_carry ));
 XOR2_X2 \stage2/gen_csa[5].FA1/HA1/_1_  (.A(ground),
    .B(sum_s1[5]),
    .Z(\stage2/gen_csa[5].FA1/ha1_sum ));
 AND2_X1 \stage2/gen_csa[5].FA1/HA2/_0_  (.A1(\stage2/gen_csa[5].FA1/ha1_sum ),
    .A2(\stage2/_07_ ),
    .ZN(\stage2/gen_csa[5].FA1/ha2_carry ));
 XOR2_X1 \stage2/gen_csa[5].FA1/HA2/_1_  (.A(\stage2/gen_csa[5].FA1/ha1_sum ),
    .B(\stage2/_07_ ),
    .Z(\stage2/sum1 [5]));
 OR2_X1 \stage2/gen_csa[5].FA1/_0_  (.A1(\stage2/gen_csa[5].FA1/ha1_carry ),
    .A2(\stage2/gen_csa[5].FA1/ha2_carry ),
    .ZN(\stage2/carry1 [5]));
 AND2_X1 \stage2/gen_csa[6].FA0/HA1/_0_  (.A1(ground),
    .A2(sum_s1[6]),
    .ZN(\stage2/gen_csa[6].FA0/ha1_carry ));
 XOR2_X2 \stage2/gen_csa[6].FA0/HA1/_1_  (.A(ground),
    .B(sum_s1[6]),
    .Z(\stage2/gen_csa[6].FA0/ha1_sum ));
 AND2_X1 \stage2/gen_csa[6].FA0/HA2/_0_  (.A1(\stage2/gen_csa[6].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\stage2/gen_csa[6].FA0/ha2_carry ));
 XOR2_X1 \stage2/gen_csa[6].FA0/HA2/_1_  (.A(\stage2/gen_csa[6].FA0/ha1_sum ),
    .B(ground),
    .Z(\stage2/sum0 [6]));
 OR2_X1 \stage2/gen_csa[6].FA0/_0_  (.A1(\stage2/gen_csa[6].FA0/ha1_carry ),
    .A2(\stage2/gen_csa[6].FA0/ha2_carry ),
    .ZN(\stage2/carry0 [6]));
 AND2_X1 \stage2/gen_csa[6].FA1/HA1/_0_  (.A1(ground),
    .A2(sum_s1[6]),
    .ZN(\stage2/gen_csa[6].FA1/ha1_carry ));
 XOR2_X2 \stage2/gen_csa[6].FA1/HA1/_1_  (.A(ground),
    .B(sum_s1[6]),
    .Z(\stage2/gen_csa[6].FA1/ha1_sum ));
 AND2_X1 \stage2/gen_csa[6].FA1/HA2/_0_  (.A1(\stage2/gen_csa[6].FA1/ha1_sum ),
    .A2(\stage2/_07_ ),
    .ZN(\stage2/gen_csa[6].FA1/ha2_carry ));
 XOR2_X1 \stage2/gen_csa[6].FA1/HA2/_1_  (.A(\stage2/gen_csa[6].FA1/ha1_sum ),
    .B(\stage2/_07_ ),
    .Z(\stage2/sum1 [6]));
 OR2_X1 \stage2/gen_csa[6].FA1/_0_  (.A1(\stage2/gen_csa[6].FA1/ha1_carry ),
    .A2(\stage2/gen_csa[6].FA1/ha2_carry ),
    .ZN(\stage2/carry1 [6]));
 AND2_X1 \stage2/gen_csa[7].FA0/HA1/_0_  (.A1(ground),
    .A2(sum_s1[7]),
    .ZN(\stage2/gen_csa[7].FA0/ha1_carry ));
 XOR2_X2 \stage2/gen_csa[7].FA0/HA1/_1_  (.A(ground),
    .B(sum_s1[7]),
    .Z(\stage2/gen_csa[7].FA0/ha1_sum ));
 AND2_X1 \stage2/gen_csa[7].FA0/HA2/_0_  (.A1(\stage2/gen_csa[7].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\stage2/gen_csa[7].FA0/ha2_carry ));
 XOR2_X1 \stage2/gen_csa[7].FA0/HA2/_1_  (.A(\stage2/gen_csa[7].FA0/ha1_sum ),
    .B(ground),
    .Z(\stage2/sum0 [7]));
 OR2_X1 \stage2/gen_csa[7].FA0/_0_  (.A1(\stage2/gen_csa[7].FA0/ha1_carry ),
    .A2(\stage2/gen_csa[7].FA0/ha2_carry ),
    .ZN(\stage2/carry0 [7]));
 AND2_X1 \stage2/gen_csa[7].FA1/HA1/_0_  (.A1(ground),
    .A2(sum_s1[7]),
    .ZN(\stage2/gen_csa[7].FA1/ha1_carry ));
 XOR2_X2 \stage2/gen_csa[7].FA1/HA1/_1_  (.A(ground),
    .B(sum_s1[7]),
    .Z(\stage2/gen_csa[7].FA1/ha1_sum ));
 AND2_X1 \stage2/gen_csa[7].FA1/HA2/_0_  (.A1(\stage2/gen_csa[7].FA1/ha1_sum ),
    .A2(\stage2/_07_ ),
    .ZN(\stage2/gen_csa[7].FA1/ha2_carry ));
 XOR2_X1 \stage2/gen_csa[7].FA1/HA2/_1_  (.A(\stage2/gen_csa[7].FA1/ha1_sum ),
    .B(\stage2/_07_ ),
    .Z(\stage2/sum1 [7]));
 OR2_X1 \stage2/gen_csa[7].FA1/_0_  (.A1(\stage2/gen_csa[7].FA1/ha1_carry ),
    .A2(\stage2/gen_csa[7].FA1/ha2_carry ),
    .ZN(\stage2/carry1 [7]));
 AND2_X1 \stage3/FA1_0/HA1/_0_  (.A1(sum_s2[4]),
    .A2(prodm3_s2[0]),
    .ZN(\stage3/FA1_0/ha1_carry ));
 XOR2_X2 \stage3/FA1_0/HA1/_1_  (.A(sum_s2[4]),
    .B(prodm3_s2[0]),
    .Z(\stage3/FA1_0/ha1_sum ));
 AND2_X1 \stage3/FA1_0/HA2/_0_  (.A1(\stage3/FA1_0/ha1_sum ),
    .A2(\stage3/_07_ ),
    .ZN(\stage3/FA1_0/ha2_carry ));
 XOR2_X1 \stage3/FA1_0/HA2/_1_  (.A(\stage3/FA1_0/ha1_sum ),
    .B(\stage3/_07_ ),
    .Z(\stage3/sum1 [0]));
 OR2_X1 \stage3/FA1_0/_0_  (.A1(\stage3/FA1_0/ha1_carry ),
    .A2(\stage3/FA1_0/ha2_carry ),
    .ZN(\stage3/carry1 [0]));
 AND2_X1 \stage3/HA0_0/_0_  (.A1(sum_s2[4]),
    .A2(prodm3_s2[0]),
    .ZN(\stage3/carry0 [0]));
 XOR2_X1 \stage3/HA0_0/_1_  (.A(sum_s2[4]),
    .B(prodm3_s2[0]),
    .Z(\stage3/sum0 [0]));
 INV_X4 \stage3/_08_  (.A(ground),
    .ZN(\stage3/_07_ ));
 MUX2_X1 \stage3/_09_  (.A(\stage3/sum0 [0]),
    .B(\stage3/sum1 [0]),
    .S(ground),
    .Z(sums3[0]));
 MUX2_X1 \stage3/_10_  (.A(\stage3/carry0 [0]),
    .B(\stage3/carry1 [0]),
    .S(ground),
    .Z(\stage3/_00_ ));
 MUX2_X1 \stage3/_11_  (.A(\stage3/sum0 [1]),
    .B(\stage3/sum1 [1]),
    .S(\stage3/_00_ ),
    .Z(sums3[1]));
 MUX2_X1 \stage3/_12_  (.A(\stage3/carry0 [1]),
    .B(\stage3/carry1 [1]),
    .S(\stage3/_00_ ),
    .Z(\stage3/_01_ ));
 MUX2_X1 \stage3/_13_  (.A(\stage3/sum0 [2]),
    .B(\stage3/sum1 [2]),
    .S(\stage3/_01_ ),
    .Z(sums3[2]));
 MUX2_X1 \stage3/_14_  (.A(\stage3/carry0 [2]),
    .B(\stage3/carry1 [2]),
    .S(\stage3/_01_ ),
    .Z(\stage3/_02_ ));
 MUX2_X1 \stage3/_15_  (.A(\stage3/sum0 [3]),
    .B(\stage3/sum1 [3]),
    .S(\stage3/_02_ ),
    .Z(sums3[3]));
 MUX2_X2 \stage3/_16_  (.A(\stage3/carry0 [3]),
    .B(\stage3/carry1 [3]),
    .S(\stage3/_02_ ),
    .Z(\stage3/_03_ ));
 MUX2_X1 \stage3/_17_  (.A(\stage3/sum0 [4]),
    .B(\stage3/sum1 [4]),
    .S(\stage3/_03_ ),
    .Z(sums3[4]));
 MUX2_X1 \stage3/_18_  (.A(\stage3/carry0 [4]),
    .B(\stage3/carry1 [4]),
    .S(\stage3/_03_ ),
    .Z(\stage3/_04_ ));
 MUX2_X1 \stage3/_19_  (.A(\stage3/sum0 [5]),
    .B(\stage3/sum1 [5]),
    .S(\stage3/_04_ ),
    .Z(sums3[5]));
 MUX2_X1 \stage3/_20_  (.A(\stage3/carry0 [5]),
    .B(\stage3/carry1 [5]),
    .S(\stage3/_04_ ),
    .Z(\stage3/_05_ ));
 MUX2_X1 \stage3/_21_  (.A(\stage3/sum0 [6]),
    .B(\stage3/sum1 [6]),
    .S(\stage3/_05_ ),
    .Z(sums3[6]));
 MUX2_X1 \stage3/_22_  (.A(\stage3/carry0 [6]),
    .B(\stage3/carry1 [6]),
    .S(\stage3/_05_ ),
    .Z(\stage3/_06_ ));
 MUX2_X1 \stage3/_23_  (.A(\stage3/sum0 [7]),
    .B(\stage3/sum1 [7]),
    .S(\stage3/_06_ ),
    .Z(sums3[7]));
 MUX2_X1 \stage3/_24_  (.A(\stage3/carry0 [7]),
    .B(\stage3/carry1 [7]),
    .S(\stage3/_06_ ),
    .Z(overflow));
 AND2_X1 \stage3/gen_csa[1].FA0/HA1/_0_  (.A1(sum_s2[5]),
    .A2(prodm3_s2[1]),
    .ZN(\stage3/gen_csa[1].FA0/ha1_carry ));
 XOR2_X2 \stage3/gen_csa[1].FA0/HA1/_1_  (.A(sum_s2[5]),
    .B(prodm3_s2[1]),
    .Z(\stage3/gen_csa[1].FA0/ha1_sum ));
 AND2_X1 \stage3/gen_csa[1].FA0/HA2/_0_  (.A1(\stage3/gen_csa[1].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\stage3/gen_csa[1].FA0/ha2_carry ));
 XOR2_X1 \stage3/gen_csa[1].FA0/HA2/_1_  (.A(\stage3/gen_csa[1].FA0/ha1_sum ),
    .B(ground),
    .Z(\stage3/sum0 [1]));
 OR2_X1 \stage3/gen_csa[1].FA0/_0_  (.A1(\stage3/gen_csa[1].FA0/ha1_carry ),
    .A2(\stage3/gen_csa[1].FA0/ha2_carry ),
    .ZN(\stage3/carry0 [1]));
 AND2_X1 \stage3/gen_csa[1].FA1/HA1/_0_  (.A1(sum_s2[5]),
    .A2(prodm3_s2[1]),
    .ZN(\stage3/gen_csa[1].FA1/ha1_carry ));
 XOR2_X2 \stage3/gen_csa[1].FA1/HA1/_1_  (.A(sum_s2[5]),
    .B(prodm3_s2[1]),
    .Z(\stage3/gen_csa[1].FA1/ha1_sum ));
 AND2_X1 \stage3/gen_csa[1].FA1/HA2/_0_  (.A1(\stage3/gen_csa[1].FA1/ha1_sum ),
    .A2(\stage3/_07_ ),
    .ZN(\stage3/gen_csa[1].FA1/ha2_carry ));
 XOR2_X1 \stage3/gen_csa[1].FA1/HA2/_1_  (.A(\stage3/gen_csa[1].FA1/ha1_sum ),
    .B(\stage3/_07_ ),
    .Z(\stage3/sum1 [1]));
 OR2_X1 \stage3/gen_csa[1].FA1/_0_  (.A1(\stage3/gen_csa[1].FA1/ha1_carry ),
    .A2(\stage3/gen_csa[1].FA1/ha2_carry ),
    .ZN(\stage3/carry1 [1]));
 AND2_X1 \stage3/gen_csa[2].FA0/HA1/_0_  (.A1(sum_s2[6]),
    .A2(prodm3_s2[2]),
    .ZN(\stage3/gen_csa[2].FA0/ha1_carry ));
 XOR2_X2 \stage3/gen_csa[2].FA0/HA1/_1_  (.A(sum_s2[6]),
    .B(prodm3_s2[2]),
    .Z(\stage3/gen_csa[2].FA0/ha1_sum ));
 AND2_X1 \stage3/gen_csa[2].FA0/HA2/_0_  (.A1(\stage3/gen_csa[2].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\stage3/gen_csa[2].FA0/ha2_carry ));
 XOR2_X1 \stage3/gen_csa[2].FA0/HA2/_1_  (.A(\stage3/gen_csa[2].FA0/ha1_sum ),
    .B(ground),
    .Z(\stage3/sum0 [2]));
 OR2_X1 \stage3/gen_csa[2].FA0/_0_  (.A1(\stage3/gen_csa[2].FA0/ha1_carry ),
    .A2(\stage3/gen_csa[2].FA0/ha2_carry ),
    .ZN(\stage3/carry0 [2]));
 AND2_X1 \stage3/gen_csa[2].FA1/HA1/_0_  (.A1(sum_s2[6]),
    .A2(prodm3_s2[2]),
    .ZN(\stage3/gen_csa[2].FA1/ha1_carry ));
 XOR2_X2 \stage3/gen_csa[2].FA1/HA1/_1_  (.A(sum_s2[6]),
    .B(prodm3_s2[2]),
    .Z(\stage3/gen_csa[2].FA1/ha1_sum ));
 AND2_X1 \stage3/gen_csa[2].FA1/HA2/_0_  (.A1(\stage3/gen_csa[2].FA1/ha1_sum ),
    .A2(\stage3/_07_ ),
    .ZN(\stage3/gen_csa[2].FA1/ha2_carry ));
 XOR2_X1 \stage3/gen_csa[2].FA1/HA2/_1_  (.A(\stage3/gen_csa[2].FA1/ha1_sum ),
    .B(\stage3/_07_ ),
    .Z(\stage3/sum1 [2]));
 OR2_X1 \stage3/gen_csa[2].FA1/_0_  (.A1(\stage3/gen_csa[2].FA1/ha1_carry ),
    .A2(\stage3/gen_csa[2].FA1/ha2_carry ),
    .ZN(\stage3/carry1 [2]));
 AND2_X1 \stage3/gen_csa[3].FA0/HA1/_0_  (.A1(sum_s2[7]),
    .A2(prodm3_s2[3]),
    .ZN(\stage3/gen_csa[3].FA0/ha1_carry ));
 XOR2_X2 \stage3/gen_csa[3].FA0/HA1/_1_  (.A(sum_s2[7]),
    .B(prodm3_s2[3]),
    .Z(\stage3/gen_csa[3].FA0/ha1_sum ));
 AND2_X1 \stage3/gen_csa[3].FA0/HA2/_0_  (.A1(\stage3/gen_csa[3].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\stage3/gen_csa[3].FA0/ha2_carry ));
 XOR2_X1 \stage3/gen_csa[3].FA0/HA2/_1_  (.A(\stage3/gen_csa[3].FA0/ha1_sum ),
    .B(ground),
    .Z(\stage3/sum0 [3]));
 OR2_X1 \stage3/gen_csa[3].FA0/_0_  (.A1(\stage3/gen_csa[3].FA0/ha1_carry ),
    .A2(\stage3/gen_csa[3].FA0/ha2_carry ),
    .ZN(\stage3/carry0 [3]));
 AND2_X1 \stage3/gen_csa[3].FA1/HA1/_0_  (.A1(sum_s2[7]),
    .A2(prodm3_s2[3]),
    .ZN(\stage3/gen_csa[3].FA1/ha1_carry ));
 XOR2_X2 \stage3/gen_csa[3].FA1/HA1/_1_  (.A(sum_s2[7]),
    .B(prodm3_s2[3]),
    .Z(\stage3/gen_csa[3].FA1/ha1_sum ));
 AND2_X1 \stage3/gen_csa[3].FA1/HA2/_0_  (.A1(\stage3/gen_csa[3].FA1/ha1_sum ),
    .A2(\stage3/_07_ ),
    .ZN(\stage3/gen_csa[3].FA1/ha2_carry ));
 XOR2_X1 \stage3/gen_csa[3].FA1/HA2/_1_  (.A(\stage3/gen_csa[3].FA1/ha1_sum ),
    .B(\stage3/_07_ ),
    .Z(\stage3/sum1 [3]));
 OR2_X1 \stage3/gen_csa[3].FA1/_0_  (.A1(\stage3/gen_csa[3].FA1/ha1_carry ),
    .A2(\stage3/gen_csa[3].FA1/ha2_carry ),
    .ZN(\stage3/carry1 [3]));
 AND2_X1 \stage3/gen_csa[4].FA0/HA1/_0_  (.A1(_000_),
    .A2(prodm3_s2[4]),
    .ZN(\stage3/gen_csa[4].FA0/ha1_carry ));
 XOR2_X2 \stage3/gen_csa[4].FA0/HA1/_1_  (.A(_000_),
    .B(prodm3_s2[4]),
    .Z(\stage3/gen_csa[4].FA0/ha1_sum ));
 AND2_X1 \stage3/gen_csa[4].FA0/HA2/_0_  (.A1(\stage3/gen_csa[4].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\stage3/gen_csa[4].FA0/ha2_carry ));
 XOR2_X1 \stage3/gen_csa[4].FA0/HA2/_1_  (.A(\stage3/gen_csa[4].FA0/ha1_sum ),
    .B(ground),
    .Z(\stage3/sum0 [4]));
 OR2_X1 \stage3/gen_csa[4].FA0/_0_  (.A1(\stage3/gen_csa[4].FA0/ha1_carry ),
    .A2(\stage3/gen_csa[4].FA0/ha2_carry ),
    .ZN(\stage3/carry0 [4]));
 AND2_X1 \stage3/gen_csa[4].FA1/HA1/_0_  (.A1(_000_),
    .A2(prodm3_s2[4]),
    .ZN(\stage3/gen_csa[4].FA1/ha1_carry ));
 XOR2_X2 \stage3/gen_csa[4].FA1/HA1/_1_  (.A(_000_),
    .B(prodm3_s2[4]),
    .Z(\stage3/gen_csa[4].FA1/ha1_sum ));
 AND2_X1 \stage3/gen_csa[4].FA1/HA2/_0_  (.A1(\stage3/gen_csa[4].FA1/ha1_sum ),
    .A2(\stage3/_07_ ),
    .ZN(\stage3/gen_csa[4].FA1/ha2_carry ));
 XOR2_X1 \stage3/gen_csa[4].FA1/HA2/_1_  (.A(\stage3/gen_csa[4].FA1/ha1_sum ),
    .B(\stage3/_07_ ),
    .Z(\stage3/sum1 [4]));
 OR2_X1 \stage3/gen_csa[4].FA1/_0_  (.A1(\stage3/gen_csa[4].FA1/ha1_carry ),
    .A2(\stage3/gen_csa[4].FA1/ha2_carry ),
    .ZN(\stage3/carry1 [4]));
 AND2_X1 \stage3/gen_csa[5].FA0/HA1/_0_  (.A1(ground),
    .A2(prodm3_s2[5]),
    .ZN(\stage3/gen_csa[5].FA0/ha1_carry ));
 XOR2_X1 \stage3/gen_csa[5].FA0/HA1/_1_  (.A(ground),
    .B(prodm3_s2[5]),
    .Z(\stage3/gen_csa[5].FA0/ha1_sum ));
 AND2_X1 \stage3/gen_csa[5].FA0/HA2/_0_  (.A1(\stage3/gen_csa[5].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\stage3/gen_csa[5].FA0/ha2_carry ));
 XOR2_X1 \stage3/gen_csa[5].FA0/HA2/_1_  (.A(\stage3/gen_csa[5].FA0/ha1_sum ),
    .B(ground),
    .Z(\stage3/sum0 [5]));
 OR2_X1 \stage3/gen_csa[5].FA0/_0_  (.A1(\stage3/gen_csa[5].FA0/ha1_carry ),
    .A2(\stage3/gen_csa[5].FA0/ha2_carry ),
    .ZN(\stage3/carry0 [5]));
 AND2_X1 \stage3/gen_csa[5].FA1/HA1/_0_  (.A1(ground),
    .A2(prodm3_s2[5]),
    .ZN(\stage3/gen_csa[5].FA1/ha1_carry ));
 XOR2_X2 \stage3/gen_csa[5].FA1/HA1/_1_  (.A(ground),
    .B(prodm3_s2[5]),
    .Z(\stage3/gen_csa[5].FA1/ha1_sum ));
 AND2_X1 \stage3/gen_csa[5].FA1/HA2/_0_  (.A1(\stage3/gen_csa[5].FA1/ha1_sum ),
    .A2(\stage3/_07_ ),
    .ZN(\stage3/gen_csa[5].FA1/ha2_carry ));
 XOR2_X1 \stage3/gen_csa[5].FA1/HA2/_1_  (.A(\stage3/gen_csa[5].FA1/ha1_sum ),
    .B(\stage3/_07_ ),
    .Z(\stage3/sum1 [5]));
 OR2_X1 \stage3/gen_csa[5].FA1/_0_  (.A1(\stage3/gen_csa[5].FA1/ha1_carry ),
    .A2(\stage3/gen_csa[5].FA1/ha2_carry ),
    .ZN(\stage3/carry1 [5]));
 AND2_X1 \stage3/gen_csa[6].FA0/HA1/_0_  (.A1(ground),
    .A2(prodm3_s2[6]),
    .ZN(\stage3/gen_csa[6].FA0/ha1_carry ));
 XOR2_X2 \stage3/gen_csa[6].FA0/HA1/_1_  (.A(ground),
    .B(prodm3_s2[6]),
    .Z(\stage3/gen_csa[6].FA0/ha1_sum ));
 AND2_X1 \stage3/gen_csa[6].FA0/HA2/_0_  (.A1(\stage3/gen_csa[6].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\stage3/gen_csa[6].FA0/ha2_carry ));
 XOR2_X1 \stage3/gen_csa[6].FA0/HA2/_1_  (.A(\stage3/gen_csa[6].FA0/ha1_sum ),
    .B(ground),
    .Z(\stage3/sum0 [6]));
 OR2_X1 \stage3/gen_csa[6].FA0/_0_  (.A1(\stage3/gen_csa[6].FA0/ha1_carry ),
    .A2(\stage3/gen_csa[6].FA0/ha2_carry ),
    .ZN(\stage3/carry0 [6]));
 AND2_X1 \stage3/gen_csa[6].FA1/HA1/_0_  (.A1(ground),
    .A2(prodm3_s2[6]),
    .ZN(\stage3/gen_csa[6].FA1/ha1_carry ));
 XOR2_X1 \stage3/gen_csa[6].FA1/HA1/_1_  (.A(ground),
    .B(prodm3_s2[6]),
    .Z(\stage3/gen_csa[6].FA1/ha1_sum ));
 AND2_X1 \stage3/gen_csa[6].FA1/HA2/_0_  (.A1(\stage3/gen_csa[6].FA1/ha1_sum ),
    .A2(\stage3/_07_ ),
    .ZN(\stage3/gen_csa[6].FA1/ha2_carry ));
 XOR2_X1 \stage3/gen_csa[6].FA1/HA2/_1_  (.A(\stage3/gen_csa[6].FA1/ha1_sum ),
    .B(\stage3/_07_ ),
    .Z(\stage3/sum1 [6]));
 OR2_X1 \stage3/gen_csa[6].FA1/_0_  (.A1(\stage3/gen_csa[6].FA1/ha1_carry ),
    .A2(\stage3/gen_csa[6].FA1/ha2_carry ),
    .ZN(\stage3/carry1 [6]));
 AND2_X1 \stage3/gen_csa[7].FA0/HA1/_0_  (.A1(ground),
    .A2(prodm3_s2[7]),
    .ZN(\stage3/gen_csa[7].FA0/ha1_carry ));
 XOR2_X2 \stage3/gen_csa[7].FA0/HA1/_1_  (.A(ground),
    .B(prodm3_s2[7]),
    .Z(\stage3/gen_csa[7].FA0/ha1_sum ));
 AND2_X1 \stage3/gen_csa[7].FA0/HA2/_0_  (.A1(\stage3/gen_csa[7].FA0/ha1_sum ),
    .A2(ground),
    .ZN(\stage3/gen_csa[7].FA0/ha2_carry ));
 XOR2_X1 \stage3/gen_csa[7].FA0/HA2/_1_  (.A(\stage3/gen_csa[7].FA0/ha1_sum ),
    .B(ground),
    .Z(\stage3/sum0 [7]));
 OR2_X1 \stage3/gen_csa[7].FA0/_0_  (.A1(\stage3/gen_csa[7].FA0/ha1_carry ),
    .A2(\stage3/gen_csa[7].FA0/ha2_carry ),
    .ZN(\stage3/carry0 [7]));
 AND2_X1 \stage3/gen_csa[7].FA1/HA1/_0_  (.A1(ground),
    .A2(prodm3_s2[7]),
    .ZN(\stage3/gen_csa[7].FA1/ha1_carry ));
 XOR2_X2 \stage3/gen_csa[7].FA1/HA1/_1_  (.A(ground),
    .B(prodm3_s2[7]),
    .Z(\stage3/gen_csa[7].FA1/ha1_sum ));
 AND2_X1 \stage3/gen_csa[7].FA1/HA2/_0_  (.A1(\stage3/gen_csa[7].FA1/ha1_sum ),
    .A2(\stage3/_07_ ),
    .ZN(\stage3/gen_csa[7].FA1/ha2_carry ));
 XOR2_X1 \stage3/gen_csa[7].FA1/HA2/_1_  (.A(\stage3/gen_csa[7].FA1/ha1_sum ),
    .B(\stage3/_07_ ),
    .Z(\stage3/sum1 [7]));
 OR2_X1 \stage3/gen_csa[7].FA1/_0_  (.A1(\stage3/gen_csa[7].FA1/ha1_carry ),
    .A2(\stage3/gen_csa[7].FA1/ha2_carry ),
    .ZN(\stage3/carry1 [7]));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_139 ();
 BUF_X4 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 BUF_X4 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_0__leaf_clk));
 BUF_X4 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_1__leaf_clk));
 BUF_X4 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_2__leaf_clk));
 BUF_X4 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_3__leaf_clk));
 BUF_X4 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_4__leaf_clk));
 BUF_X4 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_5__leaf_clk));
 BUF_X4 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_6__leaf_clk));
 BUF_X4 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_7__leaf_clk));
 INV_X4 clkload0 (.A(clknet_3_1__leaf_clk));
 INV_X8 clkload1 (.A(clknet_3_2__leaf_clk));
 INV_X4 clkload2 (.A(clknet_3_3__leaf_clk));
 INV_X4 clkload3 (.A(clknet_3_4__leaf_clk));
 INV_X2 clkload4 (.A(clknet_3_5__leaf_clk));
 INV_X4 clkload5 (.A(clknet_3_6__leaf_clk));
 INV_X8 clkload6 (.A(clknet_3_7__leaf_clk));
endmodule
